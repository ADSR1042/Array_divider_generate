module divider_32bit(
    input wire clk,
    input wire rst,
    input wire [31:0] dividend,
    input wire [31:0] divisor,
    output wire [32:0] quotient,
    output wire [32:0] remainder
);
wire c0001,c0002,c0003,c0004,c0005,c0006,c0007,c0008,c0009,c0010,c0011,c0012,c0013,c0014,c0015,c0016,c0017,c0018,c0019,c0020,c0021,c0022,c0023,c0024,c0025,c0026,c0027,c0028,c0029,c0030,c0031,c0032;
wire c0101,c0102,c0103,c0104,c0105,c0106,c0107,c0108,c0109,c0110,c0111,c0112,c0113,c0114,c0115,c0116,c0117,c0118,c0119,c0120,c0121,c0122,c0123,c0124,c0125,c0126,c0127,c0128,c0129,c0130,c0131,c0132;
wire c0201,c0202,c0203,c0204,c0205,c0206,c0207,c0208,c0209,c0210,c0211,c0212,c0213,c0214,c0215,c0216,c0217,c0218,c0219,c0220,c0221,c0222,c0223,c0224,c0225,c0226,c0227,c0228,c0229,c0230,c0231,c0232;
wire c0301,c0302,c0303,c0304,c0305,c0306,c0307,c0308,c0309,c0310,c0311,c0312,c0313,c0314,c0315,c0316,c0317,c0318,c0319,c0320,c0321,c0322,c0323,c0324,c0325,c0326,c0327,c0328,c0329,c0330,c0331,c0332;
wire c0401,c0402,c0403,c0404,c0405,c0406,c0407,c0408,c0409,c0410,c0411,c0412,c0413,c0414,c0415,c0416,c0417,c0418,c0419,c0420,c0421,c0422,c0423,c0424,c0425,c0426,c0427,c0428,c0429,c0430,c0431,c0432;
wire c0501,c0502,c0503,c0504,c0505,c0506,c0507,c0508,c0509,c0510,c0511,c0512,c0513,c0514,c0515,c0516,c0517,c0518,c0519,c0520,c0521,c0522,c0523,c0524,c0525,c0526,c0527,c0528,c0529,c0530,c0531,c0532;
wire c0601,c0602,c0603,c0604,c0605,c0606,c0607,c0608,c0609,c0610,c0611,c0612,c0613,c0614,c0615,c0616,c0617,c0618,c0619,c0620,c0621,c0622,c0623,c0624,c0625,c0626,c0627,c0628,c0629,c0630,c0631,c0632;
wire c0701,c0702,c0703,c0704,c0705,c0706,c0707,c0708,c0709,c0710,c0711,c0712,c0713,c0714,c0715,c0716,c0717,c0718,c0719,c0720,c0721,c0722,c0723,c0724,c0725,c0726,c0727,c0728,c0729,c0730,c0731,c0732;
wire c0801,c0802,c0803,c0804,c0805,c0806,c0807,c0808,c0809,c0810,c0811,c0812,c0813,c0814,c0815,c0816,c0817,c0818,c0819,c0820,c0821,c0822,c0823,c0824,c0825,c0826,c0827,c0828,c0829,c0830,c0831,c0832;
wire c0901,c0902,c0903,c0904,c0905,c0906,c0907,c0908,c0909,c0910,c0911,c0912,c0913,c0914,c0915,c0916,c0917,c0918,c0919,c0920,c0921,c0922,c0923,c0924,c0925,c0926,c0927,c0928,c0929,c0930,c0931,c0932;
wire c1001,c1002,c1003,c1004,c1005,c1006,c1007,c1008,c1009,c1010,c1011,c1012,c1013,c1014,c1015,c1016,c1017,c1018,c1019,c1020,c1021,c1022,c1023,c1024,c1025,c1026,c1027,c1028,c1029,c1030,c1031,c1032;
wire c1101,c1102,c1103,c1104,c1105,c1106,c1107,c1108,c1109,c1110,c1111,c1112,c1113,c1114,c1115,c1116,c1117,c1118,c1119,c1120,c1121,c1122,c1123,c1124,c1125,c1126,c1127,c1128,c1129,c1130,c1131,c1132;
wire c1201,c1202,c1203,c1204,c1205,c1206,c1207,c1208,c1209,c1210,c1211,c1212,c1213,c1214,c1215,c1216,c1217,c1218,c1219,c1220,c1221,c1222,c1223,c1224,c1225,c1226,c1227,c1228,c1229,c1230,c1231,c1232;
wire c1301,c1302,c1303,c1304,c1305,c1306,c1307,c1308,c1309,c1310,c1311,c1312,c1313,c1314,c1315,c1316,c1317,c1318,c1319,c1320,c1321,c1322,c1323,c1324,c1325,c1326,c1327,c1328,c1329,c1330,c1331,c1332;
wire c1401,c1402,c1403,c1404,c1405,c1406,c1407,c1408,c1409,c1410,c1411,c1412,c1413,c1414,c1415,c1416,c1417,c1418,c1419,c1420,c1421,c1422,c1423,c1424,c1425,c1426,c1427,c1428,c1429,c1430,c1431,c1432;
wire c1501,c1502,c1503,c1504,c1505,c1506,c1507,c1508,c1509,c1510,c1511,c1512,c1513,c1514,c1515,c1516,c1517,c1518,c1519,c1520,c1521,c1522,c1523,c1524,c1525,c1526,c1527,c1528,c1529,c1530,c1531,c1532;
wire c1601,c1602,c1603,c1604,c1605,c1606,c1607,c1608,c1609,c1610,c1611,c1612,c1613,c1614,c1615,c1616,c1617,c1618,c1619,c1620,c1621,c1622,c1623,c1624,c1625,c1626,c1627,c1628,c1629,c1630,c1631,c1632;
wire c1701,c1702,c1703,c1704,c1705,c1706,c1707,c1708,c1709,c1710,c1711,c1712,c1713,c1714,c1715,c1716,c1717,c1718,c1719,c1720,c1721,c1722,c1723,c1724,c1725,c1726,c1727,c1728,c1729,c1730,c1731,c1732;
wire c1801,c1802,c1803,c1804,c1805,c1806,c1807,c1808,c1809,c1810,c1811,c1812,c1813,c1814,c1815,c1816,c1817,c1818,c1819,c1820,c1821,c1822,c1823,c1824,c1825,c1826,c1827,c1828,c1829,c1830,c1831,c1832;
wire c1901,c1902,c1903,c1904,c1905,c1906,c1907,c1908,c1909,c1910,c1911,c1912,c1913,c1914,c1915,c1916,c1917,c1918,c1919,c1920,c1921,c1922,c1923,c1924,c1925,c1926,c1927,c1928,c1929,c1930,c1931,c1932;
wire c2001,c2002,c2003,c2004,c2005,c2006,c2007,c2008,c2009,c2010,c2011,c2012,c2013,c2014,c2015,c2016,c2017,c2018,c2019,c2020,c2021,c2022,c2023,c2024,c2025,c2026,c2027,c2028,c2029,c2030,c2031,c2032;
wire c2101,c2102,c2103,c2104,c2105,c2106,c2107,c2108,c2109,c2110,c2111,c2112,c2113,c2114,c2115,c2116,c2117,c2118,c2119,c2120,c2121,c2122,c2123,c2124,c2125,c2126,c2127,c2128,c2129,c2130,c2131,c2132;
wire c2201,c2202,c2203,c2204,c2205,c2206,c2207,c2208,c2209,c2210,c2211,c2212,c2213,c2214,c2215,c2216,c2217,c2218,c2219,c2220,c2221,c2222,c2223,c2224,c2225,c2226,c2227,c2228,c2229,c2230,c2231,c2232;
wire c2301,c2302,c2303,c2304,c2305,c2306,c2307,c2308,c2309,c2310,c2311,c2312,c2313,c2314,c2315,c2316,c2317,c2318,c2319,c2320,c2321,c2322,c2323,c2324,c2325,c2326,c2327,c2328,c2329,c2330,c2331,c2332;
wire c2401,c2402,c2403,c2404,c2405,c2406,c2407,c2408,c2409,c2410,c2411,c2412,c2413,c2414,c2415,c2416,c2417,c2418,c2419,c2420,c2421,c2422,c2423,c2424,c2425,c2426,c2427,c2428,c2429,c2430,c2431,c2432;
wire c2501,c2502,c2503,c2504,c2505,c2506,c2507,c2508,c2509,c2510,c2511,c2512,c2513,c2514,c2515,c2516,c2517,c2518,c2519,c2520,c2521,c2522,c2523,c2524,c2525,c2526,c2527,c2528,c2529,c2530,c2531,c2532;
wire c2601,c2602,c2603,c2604,c2605,c2606,c2607,c2608,c2609,c2610,c2611,c2612,c2613,c2614,c2615,c2616,c2617,c2618,c2619,c2620,c2621,c2622,c2623,c2624,c2625,c2626,c2627,c2628,c2629,c2630,c2631,c2632;
wire c2701,c2702,c2703,c2704,c2705,c2706,c2707,c2708,c2709,c2710,c2711,c2712,c2713,c2714,c2715,c2716,c2717,c2718,c2719,c2720,c2721,c2722,c2723,c2724,c2725,c2726,c2727,c2728,c2729,c2730,c2731,c2732;
wire c2801,c2802,c2803,c2804,c2805,c2806,c2807,c2808,c2809,c2810,c2811,c2812,c2813,c2814,c2815,c2816,c2817,c2818,c2819,c2820,c2821,c2822,c2823,c2824,c2825,c2826,c2827,c2828,c2829,c2830,c2831,c2832;
wire c2901,c2902,c2903,c2904,c2905,c2906,c2907,c2908,c2909,c2910,c2911,c2912,c2913,c2914,c2915,c2916,c2917,c2918,c2919,c2920,c2921,c2922,c2923,c2924,c2925,c2926,c2927,c2928,c2929,c2930,c2931,c2932;
wire c3001,c3002,c3003,c3004,c3005,c3006,c3007,c3008,c3009,c3010,c3011,c3012,c3013,c3014,c3015,c3016,c3017,c3018,c3019,c3020,c3021,c3022,c3023,c3024,c3025,c3026,c3027,c3028,c3029,c3030,c3031,c3032;
wire c3101,c3102,c3103,c3104,c3105,c3106,c3107,c3108,c3109,c3110,c3111,c3112,c3113,c3114,c3115,c3116,c3117,c3118,c3119,c3120,c3121,c3122,c3123,c3124,c3125,c3126,c3127,c3128,c3129,c3130,c3131,c3132;
wire c3201,c3202,c3203,c3204,c3205,c3206,c3207,c3208,c3209,c3210,c3211,c3212,c3213,c3214,c3215,c3216,c3217,c3218,c3219,c3220,c3221,c3222,c3223,c3224,c3225,c3226,c3227,c3228,c3229,c3230,c3231,c3232;
wire s0000,s0001,s0002,s0003,s0004,s0005,s0006,s0007,s0008,s0009,s0010,s0011,s0012,s0013,s0014,s0015,s0016,s0017,s0018,s0019,s0020,s0021,s0022,s0023,s0024,s0025,s0026,s0027,s0028,s0029,s0030,s0031,s0032;
wire s0100,s0101,s0102,s0103,s0104,s0105,s0106,s0107,s0108,s0109,s0110,s0111,s0112,s0113,s0114,s0115,s0116,s0117,s0118,s0119,s0120,s0121,s0122,s0123,s0124,s0125,s0126,s0127,s0128,s0129,s0130,s0131,s0132;
wire s0200,s0201,s0202,s0203,s0204,s0205,s0206,s0207,s0208,s0209,s0210,s0211,s0212,s0213,s0214,s0215,s0216,s0217,s0218,s0219,s0220,s0221,s0222,s0223,s0224,s0225,s0226,s0227,s0228,s0229,s0230,s0231,s0232;
wire s0300,s0301,s0302,s0303,s0304,s0305,s0306,s0307,s0308,s0309,s0310,s0311,s0312,s0313,s0314,s0315,s0316,s0317,s0318,s0319,s0320,s0321,s0322,s0323,s0324,s0325,s0326,s0327,s0328,s0329,s0330,s0331,s0332;
wire s0400,s0401,s0402,s0403,s0404,s0405,s0406,s0407,s0408,s0409,s0410,s0411,s0412,s0413,s0414,s0415,s0416,s0417,s0418,s0419,s0420,s0421,s0422,s0423,s0424,s0425,s0426,s0427,s0428,s0429,s0430,s0431,s0432;
wire s0500,s0501,s0502,s0503,s0504,s0505,s0506,s0507,s0508,s0509,s0510,s0511,s0512,s0513,s0514,s0515,s0516,s0517,s0518,s0519,s0520,s0521,s0522,s0523,s0524,s0525,s0526,s0527,s0528,s0529,s0530,s0531,s0532;
wire s0600,s0601,s0602,s0603,s0604,s0605,s0606,s0607,s0608,s0609,s0610,s0611,s0612,s0613,s0614,s0615,s0616,s0617,s0618,s0619,s0620,s0621,s0622,s0623,s0624,s0625,s0626,s0627,s0628,s0629,s0630,s0631,s0632;
wire s0700,s0701,s0702,s0703,s0704,s0705,s0706,s0707,s0708,s0709,s0710,s0711,s0712,s0713,s0714,s0715,s0716,s0717,s0718,s0719,s0720,s0721,s0722,s0723,s0724,s0725,s0726,s0727,s0728,s0729,s0730,s0731,s0732;
wire s0800,s0801,s0802,s0803,s0804,s0805,s0806,s0807,s0808,s0809,s0810,s0811,s0812,s0813,s0814,s0815,s0816,s0817,s0818,s0819,s0820,s0821,s0822,s0823,s0824,s0825,s0826,s0827,s0828,s0829,s0830,s0831,s0832;
wire s0900,s0901,s0902,s0903,s0904,s0905,s0906,s0907,s0908,s0909,s0910,s0911,s0912,s0913,s0914,s0915,s0916,s0917,s0918,s0919,s0920,s0921,s0922,s0923,s0924,s0925,s0926,s0927,s0928,s0929,s0930,s0931,s0932;
wire s1000,s1001,s1002,s1003,s1004,s1005,s1006,s1007,s1008,s1009,s1010,s1011,s1012,s1013,s1014,s1015,s1016,s1017,s1018,s1019,s1020,s1021,s1022,s1023,s1024,s1025,s1026,s1027,s1028,s1029,s1030,s1031,s1032;
wire s1100,s1101,s1102,s1103,s1104,s1105,s1106,s1107,s1108,s1109,s1110,s1111,s1112,s1113,s1114,s1115,s1116,s1117,s1118,s1119,s1120,s1121,s1122,s1123,s1124,s1125,s1126,s1127,s1128,s1129,s1130,s1131,s1132;
wire s1200,s1201,s1202,s1203,s1204,s1205,s1206,s1207,s1208,s1209,s1210,s1211,s1212,s1213,s1214,s1215,s1216,s1217,s1218,s1219,s1220,s1221,s1222,s1223,s1224,s1225,s1226,s1227,s1228,s1229,s1230,s1231,s1232;
wire s1300,s1301,s1302,s1303,s1304,s1305,s1306,s1307,s1308,s1309,s1310,s1311,s1312,s1313,s1314,s1315,s1316,s1317,s1318,s1319,s1320,s1321,s1322,s1323,s1324,s1325,s1326,s1327,s1328,s1329,s1330,s1331,s1332;
wire s1400,s1401,s1402,s1403,s1404,s1405,s1406,s1407,s1408,s1409,s1410,s1411,s1412,s1413,s1414,s1415,s1416,s1417,s1418,s1419,s1420,s1421,s1422,s1423,s1424,s1425,s1426,s1427,s1428,s1429,s1430,s1431,s1432;
wire s1500,s1501,s1502,s1503,s1504,s1505,s1506,s1507,s1508,s1509,s1510,s1511,s1512,s1513,s1514,s1515,s1516,s1517,s1518,s1519,s1520,s1521,s1522,s1523,s1524,s1525,s1526,s1527,s1528,s1529,s1530,s1531,s1532;
wire s1600,s1601,s1602,s1603,s1604,s1605,s1606,s1607,s1608,s1609,s1610,s1611,s1612,s1613,s1614,s1615,s1616,s1617,s1618,s1619,s1620,s1621,s1622,s1623,s1624,s1625,s1626,s1627,s1628,s1629,s1630,s1631,s1632;
wire s1700,s1701,s1702,s1703,s1704,s1705,s1706,s1707,s1708,s1709,s1710,s1711,s1712,s1713,s1714,s1715,s1716,s1717,s1718,s1719,s1720,s1721,s1722,s1723,s1724,s1725,s1726,s1727,s1728,s1729,s1730,s1731,s1732;
wire s1800,s1801,s1802,s1803,s1804,s1805,s1806,s1807,s1808,s1809,s1810,s1811,s1812,s1813,s1814,s1815,s1816,s1817,s1818,s1819,s1820,s1821,s1822,s1823,s1824,s1825,s1826,s1827,s1828,s1829,s1830,s1831,s1832;
wire s1900,s1901,s1902,s1903,s1904,s1905,s1906,s1907,s1908,s1909,s1910,s1911,s1912,s1913,s1914,s1915,s1916,s1917,s1918,s1919,s1920,s1921,s1922,s1923,s1924,s1925,s1926,s1927,s1928,s1929,s1930,s1931,s1932;
wire s2000,s2001,s2002,s2003,s2004,s2005,s2006,s2007,s2008,s2009,s2010,s2011,s2012,s2013,s2014,s2015,s2016,s2017,s2018,s2019,s2020,s2021,s2022,s2023,s2024,s2025,s2026,s2027,s2028,s2029,s2030,s2031,s2032;
wire s2100,s2101,s2102,s2103,s2104,s2105,s2106,s2107,s2108,s2109,s2110,s2111,s2112,s2113,s2114,s2115,s2116,s2117,s2118,s2119,s2120,s2121,s2122,s2123,s2124,s2125,s2126,s2127,s2128,s2129,s2130,s2131,s2132;
wire s2200,s2201,s2202,s2203,s2204,s2205,s2206,s2207,s2208,s2209,s2210,s2211,s2212,s2213,s2214,s2215,s2216,s2217,s2218,s2219,s2220,s2221,s2222,s2223,s2224,s2225,s2226,s2227,s2228,s2229,s2230,s2231,s2232;
wire s2300,s2301,s2302,s2303,s2304,s2305,s2306,s2307,s2308,s2309,s2310,s2311,s2312,s2313,s2314,s2315,s2316,s2317,s2318,s2319,s2320,s2321,s2322,s2323,s2324,s2325,s2326,s2327,s2328,s2329,s2330,s2331,s2332;
wire s2400,s2401,s2402,s2403,s2404,s2405,s2406,s2407,s2408,s2409,s2410,s2411,s2412,s2413,s2414,s2415,s2416,s2417,s2418,s2419,s2420,s2421,s2422,s2423,s2424,s2425,s2426,s2427,s2428,s2429,s2430,s2431,s2432;
wire s2500,s2501,s2502,s2503,s2504,s2505,s2506,s2507,s2508,s2509,s2510,s2511,s2512,s2513,s2514,s2515,s2516,s2517,s2518,s2519,s2520,s2521,s2522,s2523,s2524,s2525,s2526,s2527,s2528,s2529,s2530,s2531,s2532;
wire s2600,s2601,s2602,s2603,s2604,s2605,s2606,s2607,s2608,s2609,s2610,s2611,s2612,s2613,s2614,s2615,s2616,s2617,s2618,s2619,s2620,s2621,s2622,s2623,s2624,s2625,s2626,s2627,s2628,s2629,s2630,s2631,s2632;
wire s2700,s2701,s2702,s2703,s2704,s2705,s2706,s2707,s2708,s2709,s2710,s2711,s2712,s2713,s2714,s2715,s2716,s2717,s2718,s2719,s2720,s2721,s2722,s2723,s2724,s2725,s2726,s2727,s2728,s2729,s2730,s2731,s2732;
wire s2800,s2801,s2802,s2803,s2804,s2805,s2806,s2807,s2808,s2809,s2810,s2811,s2812,s2813,s2814,s2815,s2816,s2817,s2818,s2819,s2820,s2821,s2822,s2823,s2824,s2825,s2826,s2827,s2828,s2829,s2830,s2831,s2832;
wire s2900,s2901,s2902,s2903,s2904,s2905,s2906,s2907,s2908,s2909,s2910,s2911,s2912,s2913,s2914,s2915,s2916,s2917,s2918,s2919,s2920,s2921,s2922,s2923,s2924,s2925,s2926,s2927,s2928,s2929,s2930,s2931,s2932;
wire s3000,s3001,s3002,s3003,s3004,s3005,s3006,s3007,s3008,s3009,s3010,s3011,s3012,s3013,s3014,s3015,s3016,s3017,s3018,s3019,s3020,s3021,s3022,s3023,s3024,s3025,s3026,s3027,s3028,s3029,s3030,s3031,s3032;
wire s3100,s3101,s3102,s3103,s3104,s3105,s3106,s3107,s3108,s3109,s3110,s3111,s3112,s3113,s3114,s3115,s3116,s3117,s3118,s3119,s3120,s3121,s3122,s3123,s3124,s3125,s3126,s3127,s3128,s3129,s3130,s3131,s3132;
wire s3200,s3201,s3202,s3203,s3204,s3205,s3206,s3207,s3208,s3209,s3210,s3211,s3212,s3213,s3214,s3215,s3216,s3217,s3218,s3219,s3220,s3221,s3222,s3223,s3224,s3225,s3226,s3227,s3228,s3229,s3230,s3231,s3232;

reg [64:0] y;
reg [32:0] d;

addsub a0_00(y[64], d[32], c0001, 1'b1, s0000, quotient[32]);
addsub a0_01(y[63], d[31], c0002, 1'b1, s0001, c0001);
addsub a0_02(y[62], d[30], c0003, 1'b1, s0002, c0002);
addsub a0_03(y[61], d[29], c0004, 1'b1, s0003, c0003);
addsub a0_04(y[60], d[28], c0005, 1'b1, s0004, c0004);
addsub a0_05(y[59], d[27], c0006, 1'b1, s0005, c0005);
addsub a0_06(y[58], d[26], c0007, 1'b1, s0006, c0006);
addsub a0_07(y[57], d[25], c0008, 1'b1, s0007, c0007);
addsub a0_08(y[56], d[24], c0009, 1'b1, s0008, c0008);
addsub a0_09(y[55], d[23], c0010, 1'b1, s0009, c0009);
addsub a0_10(y[54], d[22], c0011, 1'b1, s0010, c0010);
addsub a0_11(y[53], d[21], c0012, 1'b1, s0011, c0011);
addsub a0_12(y[52], d[20], c0013, 1'b1, s0012, c0012);
addsub a0_13(y[51], d[19], c0014, 1'b1, s0013, c0013);
addsub a0_14(y[50], d[18], c0015, 1'b1, s0014, c0014);
addsub a0_15(y[49], d[17], c0016, 1'b1, s0015, c0015);
addsub a0_16(y[48], d[16], c0017, 1'b1, s0016, c0016);
addsub a0_17(y[47], d[15], c0018, 1'b1, s0017, c0017);
addsub a0_18(y[46], d[14], c0019, 1'b1, s0018, c0018);
addsub a0_19(y[45], d[13], c0020, 1'b1, s0019, c0019);
addsub a0_20(y[44], d[12], c0021, 1'b1, s0020, c0020);
addsub a0_21(y[43], d[11], c0022, 1'b1, s0021, c0021);
addsub a0_22(y[42], d[10], c0023, 1'b1, s0022, c0022);
addsub a0_23(y[41], d[09], c0024, 1'b1, s0023, c0023);
addsub a0_24(y[40], d[08], c0025, 1'b1, s0024, c0024);
addsub a0_25(y[39], d[07], c0026, 1'b1, s0025, c0025);
addsub a0_26(y[38], d[06], c0027, 1'b1, s0026, c0026);
addsub a0_27(y[37], d[05], c0028, 1'b1, s0027, c0027);
addsub a0_28(y[36], d[04], c0029, 1'b1, s0028, c0028);
addsub a0_29(y[35], d[03], c0030, 1'b1, s0029, c0029);
addsub a0_30(y[34], d[02], c0031, 1'b1, s0030, c0030);
addsub a0_31(y[33], d[01], c0032, 1'b1, s0031, c0031);
addsub a0_32(y[32], d[00], 1'b1, 1'b1, s0032, c0032);


addsub a01_00(s0001, d[32], c0101, quotient[32], s0100, quotient[31]);
addsub a01_01(s0002, d[31], c0102, quotient[32], s0101, c0101);
addsub a01_02(s0003, d[30], c0103, quotient[32], s0102, c0102);
addsub a01_03(s0004, d[29], c0104, quotient[32], s0103, c0103);
addsub a01_04(s0005, d[28], c0105, quotient[32], s0104, c0104);
addsub a01_05(s0006, d[27], c0106, quotient[32], s0105, c0105);
addsub a01_06(s0007, d[26], c0107, quotient[32], s0106, c0106);
addsub a01_07(s0008, d[25], c0108, quotient[32], s0107, c0107);
addsub a01_08(s0009, d[24], c0109, quotient[32], s0108, c0108);
addsub a01_09(s0010, d[23], c0110, quotient[32], s0109, c0109);
addsub a01_10(s0011, d[22], c0111, quotient[32], s0110, c0110);
addsub a01_11(s0012, d[21], c0112, quotient[32], s0111, c0111);
addsub a01_12(s0013, d[20], c0113, quotient[32], s0112, c0112);
addsub a01_13(s0014, d[19], c0114, quotient[32], s0113, c0113);
addsub a01_14(s0015, d[18], c0115, quotient[32], s0114, c0114);
addsub a01_15(s0016, d[17], c0116, quotient[32], s0115, c0115);
addsub a01_16(s0017, d[16], c0117, quotient[32], s0116, c0116);
addsub a01_17(s0018, d[15], c0118, quotient[32], s0117, c0117);
addsub a01_18(s0019, d[14], c0119, quotient[32], s0118, c0118);
addsub a01_19(s0020, d[13], c0120, quotient[32], s0119, c0119);
addsub a01_20(s0021, d[12], c0121, quotient[32], s0120, c0120);
addsub a01_21(s0022, d[11], c0122, quotient[32], s0121, c0121);
addsub a01_22(s0023, d[10], c0123, quotient[32], s0122, c0122);
addsub a01_23(s0024, d[09], c0124, quotient[32], s0123, c0123);
addsub a01_24(s0025, d[08], c0125, quotient[32], s0124, c0124);
addsub a01_25(s0026, d[07], c0126, quotient[32], s0125, c0125);
addsub a01_26(s0027, d[06], c0127, quotient[32], s0126, c0126);
addsub a01_27(s0028, d[05], c0128, quotient[32], s0127, c0127);
addsub a01_28(s0029, d[04], c0129, quotient[32], s0128, c0128);
addsub a01_29(s0030, d[03], c0130, quotient[32], s0129, c0129);
addsub a01_30(s0031, d[02], c0131, quotient[32], s0130, c0130);
addsub a01_31(s0032, d[01], c0132, quotient[32], s0131, c0131);
addsub a01_32(y[31], d[00], quotient[32], quotient[32], s0132, c0132);


addsub a02_00(s0101, d[32], c0201, quotient[31], s0200, quotient[30]);
addsub a02_01(s0102, d[31], c0202, quotient[31], s0201, c0201);
addsub a02_02(s0103, d[30], c0203, quotient[31], s0202, c0202);
addsub a02_03(s0104, d[29], c0204, quotient[31], s0203, c0203);
addsub a02_04(s0105, d[28], c0205, quotient[31], s0204, c0204);
addsub a02_05(s0106, d[27], c0206, quotient[31], s0205, c0205);
addsub a02_06(s0107, d[26], c0207, quotient[31], s0206, c0206);
addsub a02_07(s0108, d[25], c0208, quotient[31], s0207, c0207);
addsub a02_08(s0109, d[24], c0209, quotient[31], s0208, c0208);
addsub a02_09(s0110, d[23], c0210, quotient[31], s0209, c0209);
addsub a02_10(s0111, d[22], c0211, quotient[31], s0210, c0210);
addsub a02_11(s0112, d[21], c0212, quotient[31], s0211, c0211);
addsub a02_12(s0113, d[20], c0213, quotient[31], s0212, c0212);
addsub a02_13(s0114, d[19], c0214, quotient[31], s0213, c0213);
addsub a02_14(s0115, d[18], c0215, quotient[31], s0214, c0214);
addsub a02_15(s0116, d[17], c0216, quotient[31], s0215, c0215);
addsub a02_16(s0117, d[16], c0217, quotient[31], s0216, c0216);
addsub a02_17(s0118, d[15], c0218, quotient[31], s0217, c0217);
addsub a02_18(s0119, d[14], c0219, quotient[31], s0218, c0218);
addsub a02_19(s0120, d[13], c0220, quotient[31], s0219, c0219);
addsub a02_20(s0121, d[12], c0221, quotient[31], s0220, c0220);
addsub a02_21(s0122, d[11], c0222, quotient[31], s0221, c0221);
addsub a02_22(s0123, d[10], c0223, quotient[31], s0222, c0222);
addsub a02_23(s0124, d[09], c0224, quotient[31], s0223, c0223);
addsub a02_24(s0125, d[08], c0225, quotient[31], s0224, c0224);
addsub a02_25(s0126, d[07], c0226, quotient[31], s0225, c0225);
addsub a02_26(s0127, d[06], c0227, quotient[31], s0226, c0226);
addsub a02_27(s0128, d[05], c0228, quotient[31], s0227, c0227);
addsub a02_28(s0129, d[04], c0229, quotient[31], s0228, c0228);
addsub a02_29(s0130, d[03], c0230, quotient[31], s0229, c0229);
addsub a02_30(s0131, d[02], c0231, quotient[31], s0230, c0230);
addsub a02_31(s0132, d[01], c0232, quotient[31], s0231, c0231);
addsub a02_32(y[30], d[00], quotient[31], quotient[31], s0232, c0232);


addsub a03_00(s0201, d[32], c0301, quotient[30], s0300, quotient[29]);
addsub a03_01(s0202, d[31], c0302, quotient[30], s0301, c0301);
addsub a03_02(s0203, d[30], c0303, quotient[30], s0302, c0302);
addsub a03_03(s0204, d[29], c0304, quotient[30], s0303, c0303);
addsub a03_04(s0205, d[28], c0305, quotient[30], s0304, c0304);
addsub a03_05(s0206, d[27], c0306, quotient[30], s0305, c0305);
addsub a03_06(s0207, d[26], c0307, quotient[30], s0306, c0306);
addsub a03_07(s0208, d[25], c0308, quotient[30], s0307, c0307);
addsub a03_08(s0209, d[24], c0309, quotient[30], s0308, c0308);
addsub a03_09(s0210, d[23], c0310, quotient[30], s0309, c0309);
addsub a03_10(s0211, d[22], c0311, quotient[30], s0310, c0310);
addsub a03_11(s0212, d[21], c0312, quotient[30], s0311, c0311);
addsub a03_12(s0213, d[20], c0313, quotient[30], s0312, c0312);
addsub a03_13(s0214, d[19], c0314, quotient[30], s0313, c0313);
addsub a03_14(s0215, d[18], c0315, quotient[30], s0314, c0314);
addsub a03_15(s0216, d[17], c0316, quotient[30], s0315, c0315);
addsub a03_16(s0217, d[16], c0317, quotient[30], s0316, c0316);
addsub a03_17(s0218, d[15], c0318, quotient[30], s0317, c0317);
addsub a03_18(s0219, d[14], c0319, quotient[30], s0318, c0318);
addsub a03_19(s0220, d[13], c0320, quotient[30], s0319, c0319);
addsub a03_20(s0221, d[12], c0321, quotient[30], s0320, c0320);
addsub a03_21(s0222, d[11], c0322, quotient[30], s0321, c0321);
addsub a03_22(s0223, d[10], c0323, quotient[30], s0322, c0322);
addsub a03_23(s0224, d[09], c0324, quotient[30], s0323, c0323);
addsub a03_24(s0225, d[08], c0325, quotient[30], s0324, c0324);
addsub a03_25(s0226, d[07], c0326, quotient[30], s0325, c0325);
addsub a03_26(s0227, d[06], c0327, quotient[30], s0326, c0326);
addsub a03_27(s0228, d[05], c0328, quotient[30], s0327, c0327);
addsub a03_28(s0229, d[04], c0329, quotient[30], s0328, c0328);
addsub a03_29(s0230, d[03], c0330, quotient[30], s0329, c0329);
addsub a03_30(s0231, d[02], c0331, quotient[30], s0330, c0330);
addsub a03_31(s0232, d[01], c0332, quotient[30], s0331, c0331);
addsub a03_32(y[29], d[00], quotient[30], quotient[30], s0332, c0332);


addsub a04_00(s0301, d[32], c0401, quotient[29], s0400, quotient[28]);
addsub a04_01(s0302, d[31], c0402, quotient[29], s0401, c0401);
addsub a04_02(s0303, d[30], c0403, quotient[29], s0402, c0402);
addsub a04_03(s0304, d[29], c0404, quotient[29], s0403, c0403);
addsub a04_04(s0305, d[28], c0405, quotient[29], s0404, c0404);
addsub a04_05(s0306, d[27], c0406, quotient[29], s0405, c0405);
addsub a04_06(s0307, d[26], c0407, quotient[29], s0406, c0406);
addsub a04_07(s0308, d[25], c0408, quotient[29], s0407, c0407);
addsub a04_08(s0309, d[24], c0409, quotient[29], s0408, c0408);
addsub a04_09(s0310, d[23], c0410, quotient[29], s0409, c0409);
addsub a04_10(s0311, d[22], c0411, quotient[29], s0410, c0410);
addsub a04_11(s0312, d[21], c0412, quotient[29], s0411, c0411);
addsub a04_12(s0313, d[20], c0413, quotient[29], s0412, c0412);
addsub a04_13(s0314, d[19], c0414, quotient[29], s0413, c0413);
addsub a04_14(s0315, d[18], c0415, quotient[29], s0414, c0414);
addsub a04_15(s0316, d[17], c0416, quotient[29], s0415, c0415);
addsub a04_16(s0317, d[16], c0417, quotient[29], s0416, c0416);
addsub a04_17(s0318, d[15], c0418, quotient[29], s0417, c0417);
addsub a04_18(s0319, d[14], c0419, quotient[29], s0418, c0418);
addsub a04_19(s0320, d[13], c0420, quotient[29], s0419, c0419);
addsub a04_20(s0321, d[12], c0421, quotient[29], s0420, c0420);
addsub a04_21(s0322, d[11], c0422, quotient[29], s0421, c0421);
addsub a04_22(s0323, d[10], c0423, quotient[29], s0422, c0422);
addsub a04_23(s0324, d[09], c0424, quotient[29], s0423, c0423);
addsub a04_24(s0325, d[08], c0425, quotient[29], s0424, c0424);
addsub a04_25(s0326, d[07], c0426, quotient[29], s0425, c0425);
addsub a04_26(s0327, d[06], c0427, quotient[29], s0426, c0426);
addsub a04_27(s0328, d[05], c0428, quotient[29], s0427, c0427);
addsub a04_28(s0329, d[04], c0429, quotient[29], s0428, c0428);
addsub a04_29(s0330, d[03], c0430, quotient[29], s0429, c0429);
addsub a04_30(s0331, d[02], c0431, quotient[29], s0430, c0430);
addsub a04_31(s0332, d[01], c0432, quotient[29], s0431, c0431);
addsub a04_32(y[28], d[00], quotient[29], quotient[29], s0432, c0432);


addsub a05_00(s0401, d[32], c0501, quotient[28], s0500, quotient[27]);
addsub a05_01(s0402, d[31], c0502, quotient[28], s0501, c0501);
addsub a05_02(s0403, d[30], c0503, quotient[28], s0502, c0502);
addsub a05_03(s0404, d[29], c0504, quotient[28], s0503, c0503);
addsub a05_04(s0405, d[28], c0505, quotient[28], s0504, c0504);
addsub a05_05(s0406, d[27], c0506, quotient[28], s0505, c0505);
addsub a05_06(s0407, d[26], c0507, quotient[28], s0506, c0506);
addsub a05_07(s0408, d[25], c0508, quotient[28], s0507, c0507);
addsub a05_08(s0409, d[24], c0509, quotient[28], s0508, c0508);
addsub a05_09(s0410, d[23], c0510, quotient[28], s0509, c0509);
addsub a05_10(s0411, d[22], c0511, quotient[28], s0510, c0510);
addsub a05_11(s0412, d[21], c0512, quotient[28], s0511, c0511);
addsub a05_12(s0413, d[20], c0513, quotient[28], s0512, c0512);
addsub a05_13(s0414, d[19], c0514, quotient[28], s0513, c0513);
addsub a05_14(s0415, d[18], c0515, quotient[28], s0514, c0514);
addsub a05_15(s0416, d[17], c0516, quotient[28], s0515, c0515);
addsub a05_16(s0417, d[16], c0517, quotient[28], s0516, c0516);
addsub a05_17(s0418, d[15], c0518, quotient[28], s0517, c0517);
addsub a05_18(s0419, d[14], c0519, quotient[28], s0518, c0518);
addsub a05_19(s0420, d[13], c0520, quotient[28], s0519, c0519);
addsub a05_20(s0421, d[12], c0521, quotient[28], s0520, c0520);
addsub a05_21(s0422, d[11], c0522, quotient[28], s0521, c0521);
addsub a05_22(s0423, d[10], c0523, quotient[28], s0522, c0522);
addsub a05_23(s0424, d[09], c0524, quotient[28], s0523, c0523);
addsub a05_24(s0425, d[08], c0525, quotient[28], s0524, c0524);
addsub a05_25(s0426, d[07], c0526, quotient[28], s0525, c0525);
addsub a05_26(s0427, d[06], c0527, quotient[28], s0526, c0526);
addsub a05_27(s0428, d[05], c0528, quotient[28], s0527, c0527);
addsub a05_28(s0429, d[04], c0529, quotient[28], s0528, c0528);
addsub a05_29(s0430, d[03], c0530, quotient[28], s0529, c0529);
addsub a05_30(s0431, d[02], c0531, quotient[28], s0530, c0530);
addsub a05_31(s0432, d[01], c0532, quotient[28], s0531, c0531);
addsub a05_32(y[27], d[00], quotient[28], quotient[28], s0532, c0532);


addsub a06_00(s0501, d[32], c0601, quotient[27], s0600, quotient[26]);
addsub a06_01(s0502, d[31], c0602, quotient[27], s0601, c0601);
addsub a06_02(s0503, d[30], c0603, quotient[27], s0602, c0602);
addsub a06_03(s0504, d[29], c0604, quotient[27], s0603, c0603);
addsub a06_04(s0505, d[28], c0605, quotient[27], s0604, c0604);
addsub a06_05(s0506, d[27], c0606, quotient[27], s0605, c0605);
addsub a06_06(s0507, d[26], c0607, quotient[27], s0606, c0606);
addsub a06_07(s0508, d[25], c0608, quotient[27], s0607, c0607);
addsub a06_08(s0509, d[24], c0609, quotient[27], s0608, c0608);
addsub a06_09(s0510, d[23], c0610, quotient[27], s0609, c0609);
addsub a06_10(s0511, d[22], c0611, quotient[27], s0610, c0610);
addsub a06_11(s0512, d[21], c0612, quotient[27], s0611, c0611);
addsub a06_12(s0513, d[20], c0613, quotient[27], s0612, c0612);
addsub a06_13(s0514, d[19], c0614, quotient[27], s0613, c0613);
addsub a06_14(s0515, d[18], c0615, quotient[27], s0614, c0614);
addsub a06_15(s0516, d[17], c0616, quotient[27], s0615, c0615);
addsub a06_16(s0517, d[16], c0617, quotient[27], s0616, c0616);
addsub a06_17(s0518, d[15], c0618, quotient[27], s0617, c0617);
addsub a06_18(s0519, d[14], c0619, quotient[27], s0618, c0618);
addsub a06_19(s0520, d[13], c0620, quotient[27], s0619, c0619);
addsub a06_20(s0521, d[12], c0621, quotient[27], s0620, c0620);
addsub a06_21(s0522, d[11], c0622, quotient[27], s0621, c0621);
addsub a06_22(s0523, d[10], c0623, quotient[27], s0622, c0622);
addsub a06_23(s0524, d[09], c0624, quotient[27], s0623, c0623);
addsub a06_24(s0525, d[08], c0625, quotient[27], s0624, c0624);
addsub a06_25(s0526, d[07], c0626, quotient[27], s0625, c0625);
addsub a06_26(s0527, d[06], c0627, quotient[27], s0626, c0626);
addsub a06_27(s0528, d[05], c0628, quotient[27], s0627, c0627);
addsub a06_28(s0529, d[04], c0629, quotient[27], s0628, c0628);
addsub a06_29(s0530, d[03], c0630, quotient[27], s0629, c0629);
addsub a06_30(s0531, d[02], c0631, quotient[27], s0630, c0630);
addsub a06_31(s0532, d[01], c0632, quotient[27], s0631, c0631);
addsub a06_32(y[26], d[00], quotient[27], quotient[27], s0632, c0632);


addsub a07_00(s0601, d[32], c0701, quotient[26], s0700, quotient[25]);
addsub a07_01(s0602, d[31], c0702, quotient[26], s0701, c0701);
addsub a07_02(s0603, d[30], c0703, quotient[26], s0702, c0702);
addsub a07_03(s0604, d[29], c0704, quotient[26], s0703, c0703);
addsub a07_04(s0605, d[28], c0705, quotient[26], s0704, c0704);
addsub a07_05(s0606, d[27], c0706, quotient[26], s0705, c0705);
addsub a07_06(s0607, d[26], c0707, quotient[26], s0706, c0706);
addsub a07_07(s0608, d[25], c0708, quotient[26], s0707, c0707);
addsub a07_08(s0609, d[24], c0709, quotient[26], s0708, c0708);
addsub a07_09(s0610, d[23], c0710, quotient[26], s0709, c0709);
addsub a07_10(s0611, d[22], c0711, quotient[26], s0710, c0710);
addsub a07_11(s0612, d[21], c0712, quotient[26], s0711, c0711);
addsub a07_12(s0613, d[20], c0713, quotient[26], s0712, c0712);
addsub a07_13(s0614, d[19], c0714, quotient[26], s0713, c0713);
addsub a07_14(s0615, d[18], c0715, quotient[26], s0714, c0714);
addsub a07_15(s0616, d[17], c0716, quotient[26], s0715, c0715);
addsub a07_16(s0617, d[16], c0717, quotient[26], s0716, c0716);
addsub a07_17(s0618, d[15], c0718, quotient[26], s0717, c0717);
addsub a07_18(s0619, d[14], c0719, quotient[26], s0718, c0718);
addsub a07_19(s0620, d[13], c0720, quotient[26], s0719, c0719);
addsub a07_20(s0621, d[12], c0721, quotient[26], s0720, c0720);
addsub a07_21(s0622, d[11], c0722, quotient[26], s0721, c0721);
addsub a07_22(s0623, d[10], c0723, quotient[26], s0722, c0722);
addsub a07_23(s0624, d[09], c0724, quotient[26], s0723, c0723);
addsub a07_24(s0625, d[08], c0725, quotient[26], s0724, c0724);
addsub a07_25(s0626, d[07], c0726, quotient[26], s0725, c0725);
addsub a07_26(s0627, d[06], c0727, quotient[26], s0726, c0726);
addsub a07_27(s0628, d[05], c0728, quotient[26], s0727, c0727);
addsub a07_28(s0629, d[04], c0729, quotient[26], s0728, c0728);
addsub a07_29(s0630, d[03], c0730, quotient[26], s0729, c0729);
addsub a07_30(s0631, d[02], c0731, quotient[26], s0730, c0730);
addsub a07_31(s0632, d[01], c0732, quotient[26], s0731, c0731);
addsub a07_32(y[25], d[00], quotient[26], quotient[26], s0732, c0732);


addsub a08_00(s0701, d[32], c0801, quotient[25], s0800, quotient[24]);
addsub a08_01(s0702, d[31], c0802, quotient[25], s0801, c0801);
addsub a08_02(s0703, d[30], c0803, quotient[25], s0802, c0802);
addsub a08_03(s0704, d[29], c0804, quotient[25], s0803, c0803);
addsub a08_04(s0705, d[28], c0805, quotient[25], s0804, c0804);
addsub a08_05(s0706, d[27], c0806, quotient[25], s0805, c0805);
addsub a08_06(s0707, d[26], c0807, quotient[25], s0806, c0806);
addsub a08_07(s0708, d[25], c0808, quotient[25], s0807, c0807);
addsub a08_08(s0709, d[24], c0809, quotient[25], s0808, c0808);
addsub a08_09(s0710, d[23], c0810, quotient[25], s0809, c0809);
addsub a08_10(s0711, d[22], c0811, quotient[25], s0810, c0810);
addsub a08_11(s0712, d[21], c0812, quotient[25], s0811, c0811);
addsub a08_12(s0713, d[20], c0813, quotient[25], s0812, c0812);
addsub a08_13(s0714, d[19], c0814, quotient[25], s0813, c0813);
addsub a08_14(s0715, d[18], c0815, quotient[25], s0814, c0814);
addsub a08_15(s0716, d[17], c0816, quotient[25], s0815, c0815);
addsub a08_16(s0717, d[16], c0817, quotient[25], s0816, c0816);
addsub a08_17(s0718, d[15], c0818, quotient[25], s0817, c0817);
addsub a08_18(s0719, d[14], c0819, quotient[25], s0818, c0818);
addsub a08_19(s0720, d[13], c0820, quotient[25], s0819, c0819);
addsub a08_20(s0721, d[12], c0821, quotient[25], s0820, c0820);
addsub a08_21(s0722, d[11], c0822, quotient[25], s0821, c0821);
addsub a08_22(s0723, d[10], c0823, quotient[25], s0822, c0822);
addsub a08_23(s0724, d[09], c0824, quotient[25], s0823, c0823);
addsub a08_24(s0725, d[08], c0825, quotient[25], s0824, c0824);
addsub a08_25(s0726, d[07], c0826, quotient[25], s0825, c0825);
addsub a08_26(s0727, d[06], c0827, quotient[25], s0826, c0826);
addsub a08_27(s0728, d[05], c0828, quotient[25], s0827, c0827);
addsub a08_28(s0729, d[04], c0829, quotient[25], s0828, c0828);
addsub a08_29(s0730, d[03], c0830, quotient[25], s0829, c0829);
addsub a08_30(s0731, d[02], c0831, quotient[25], s0830, c0830);
addsub a08_31(s0732, d[01], c0832, quotient[25], s0831, c0831);
addsub a08_32(y[24], d[00], quotient[25], quotient[25], s0832, c0832);


addsub a09_00(s0801, d[32], c0901, quotient[24], s0900, quotient[23]);
addsub a09_01(s0802, d[31], c0902, quotient[24], s0901, c0901);
addsub a09_02(s0803, d[30], c0903, quotient[24], s0902, c0902);
addsub a09_03(s0804, d[29], c0904, quotient[24], s0903, c0903);
addsub a09_04(s0805, d[28], c0905, quotient[24], s0904, c0904);
addsub a09_05(s0806, d[27], c0906, quotient[24], s0905, c0905);
addsub a09_06(s0807, d[26], c0907, quotient[24], s0906, c0906);
addsub a09_07(s0808, d[25], c0908, quotient[24], s0907, c0907);
addsub a09_08(s0809, d[24], c0909, quotient[24], s0908, c0908);
addsub a09_09(s0810, d[23], c0910, quotient[24], s0909, c0909);
addsub a09_10(s0811, d[22], c0911, quotient[24], s0910, c0910);
addsub a09_11(s0812, d[21], c0912, quotient[24], s0911, c0911);
addsub a09_12(s0813, d[20], c0913, quotient[24], s0912, c0912);
addsub a09_13(s0814, d[19], c0914, quotient[24], s0913, c0913);
addsub a09_14(s0815, d[18], c0915, quotient[24], s0914, c0914);
addsub a09_15(s0816, d[17], c0916, quotient[24], s0915, c0915);
addsub a09_16(s0817, d[16], c0917, quotient[24], s0916, c0916);
addsub a09_17(s0818, d[15], c0918, quotient[24], s0917, c0917);
addsub a09_18(s0819, d[14], c0919, quotient[24], s0918, c0918);
addsub a09_19(s0820, d[13], c0920, quotient[24], s0919, c0919);
addsub a09_20(s0821, d[12], c0921, quotient[24], s0920, c0920);
addsub a09_21(s0822, d[11], c0922, quotient[24], s0921, c0921);
addsub a09_22(s0823, d[10], c0923, quotient[24], s0922, c0922);
addsub a09_23(s0824, d[09], c0924, quotient[24], s0923, c0923);
addsub a09_24(s0825, d[08], c0925, quotient[24], s0924, c0924);
addsub a09_25(s0826, d[07], c0926, quotient[24], s0925, c0925);
addsub a09_26(s0827, d[06], c0927, quotient[24], s0926, c0926);
addsub a09_27(s0828, d[05], c0928, quotient[24], s0927, c0927);
addsub a09_28(s0829, d[04], c0929, quotient[24], s0928, c0928);
addsub a09_29(s0830, d[03], c0930, quotient[24], s0929, c0929);
addsub a09_30(s0831, d[02], c0931, quotient[24], s0930, c0930);
addsub a09_31(s0832, d[01], c0932, quotient[24], s0931, c0931);
addsub a09_32(y[23], d[00], quotient[24], quotient[24], s0932, c0932);


addsub a10_00(s0901, d[32], c1001, quotient[23], s1000, quotient[22]);
addsub a10_01(s0902, d[31], c1002, quotient[23], s1001, c1001);
addsub a10_02(s0903, d[30], c1003, quotient[23], s1002, c1002);
addsub a10_03(s0904, d[29], c1004, quotient[23], s1003, c1003);
addsub a10_04(s0905, d[28], c1005, quotient[23], s1004, c1004);
addsub a10_05(s0906, d[27], c1006, quotient[23], s1005, c1005);
addsub a10_06(s0907, d[26], c1007, quotient[23], s1006, c1006);
addsub a10_07(s0908, d[25], c1008, quotient[23], s1007, c1007);
addsub a10_08(s0909, d[24], c1009, quotient[23], s1008, c1008);
addsub a10_09(s0910, d[23], c1010, quotient[23], s1009, c1009);
addsub a10_10(s0911, d[22], c1011, quotient[23], s1010, c1010);
addsub a10_11(s0912, d[21], c1012, quotient[23], s1011, c1011);
addsub a10_12(s0913, d[20], c1013, quotient[23], s1012, c1012);
addsub a10_13(s0914, d[19], c1014, quotient[23], s1013, c1013);
addsub a10_14(s0915, d[18], c1015, quotient[23], s1014, c1014);
addsub a10_15(s0916, d[17], c1016, quotient[23], s1015, c1015);
addsub a10_16(s0917, d[16], c1017, quotient[23], s1016, c1016);
addsub a10_17(s0918, d[15], c1018, quotient[23], s1017, c1017);
addsub a10_18(s0919, d[14], c1019, quotient[23], s1018, c1018);
addsub a10_19(s0920, d[13], c1020, quotient[23], s1019, c1019);
addsub a10_20(s0921, d[12], c1021, quotient[23], s1020, c1020);
addsub a10_21(s0922, d[11], c1022, quotient[23], s1021, c1021);
addsub a10_22(s0923, d[10], c1023, quotient[23], s1022, c1022);
addsub a10_23(s0924, d[09], c1024, quotient[23], s1023, c1023);
addsub a10_24(s0925, d[08], c1025, quotient[23], s1024, c1024);
addsub a10_25(s0926, d[07], c1026, quotient[23], s1025, c1025);
addsub a10_26(s0927, d[06], c1027, quotient[23], s1026, c1026);
addsub a10_27(s0928, d[05], c1028, quotient[23], s1027, c1027);
addsub a10_28(s0929, d[04], c1029, quotient[23], s1028, c1028);
addsub a10_29(s0930, d[03], c1030, quotient[23], s1029, c1029);
addsub a10_30(s0931, d[02], c1031, quotient[23], s1030, c1030);
addsub a10_31(s0932, d[01], c1032, quotient[23], s1031, c1031);
addsub a10_32(y[22], d[00], quotient[23], quotient[23], s1032, c1032);


addsub a11_00(s1001, d[32], c1101, quotient[22], s1100, quotient[21]);
addsub a11_01(s1002, d[31], c1102, quotient[22], s1101, c1101);
addsub a11_02(s1003, d[30], c1103, quotient[22], s1102, c1102);
addsub a11_03(s1004, d[29], c1104, quotient[22], s1103, c1103);
addsub a11_04(s1005, d[28], c1105, quotient[22], s1104, c1104);
addsub a11_05(s1006, d[27], c1106, quotient[22], s1105, c1105);
addsub a11_06(s1007, d[26], c1107, quotient[22], s1106, c1106);
addsub a11_07(s1008, d[25], c1108, quotient[22], s1107, c1107);
addsub a11_08(s1009, d[24], c1109, quotient[22], s1108, c1108);
addsub a11_09(s1010, d[23], c1110, quotient[22], s1109, c1109);
addsub a11_10(s1011, d[22], c1111, quotient[22], s1110, c1110);
addsub a11_11(s1012, d[21], c1112, quotient[22], s1111, c1111);
addsub a11_12(s1013, d[20], c1113, quotient[22], s1112, c1112);
addsub a11_13(s1014, d[19], c1114, quotient[22], s1113, c1113);
addsub a11_14(s1015, d[18], c1115, quotient[22], s1114, c1114);
addsub a11_15(s1016, d[17], c1116, quotient[22], s1115, c1115);
addsub a11_16(s1017, d[16], c1117, quotient[22], s1116, c1116);
addsub a11_17(s1018, d[15], c1118, quotient[22], s1117, c1117);
addsub a11_18(s1019, d[14], c1119, quotient[22], s1118, c1118);
addsub a11_19(s1020, d[13], c1120, quotient[22], s1119, c1119);
addsub a11_20(s1021, d[12], c1121, quotient[22], s1120, c1120);
addsub a11_21(s1022, d[11], c1122, quotient[22], s1121, c1121);
addsub a11_22(s1023, d[10], c1123, quotient[22], s1122, c1122);
addsub a11_23(s1024, d[09], c1124, quotient[22], s1123, c1123);
addsub a11_24(s1025, d[08], c1125, quotient[22], s1124, c1124);
addsub a11_25(s1026, d[07], c1126, quotient[22], s1125, c1125);
addsub a11_26(s1027, d[06], c1127, quotient[22], s1126, c1126);
addsub a11_27(s1028, d[05], c1128, quotient[22], s1127, c1127);
addsub a11_28(s1029, d[04], c1129, quotient[22], s1128, c1128);
addsub a11_29(s1030, d[03], c1130, quotient[22], s1129, c1129);
addsub a11_30(s1031, d[02], c1131, quotient[22], s1130, c1130);
addsub a11_31(s1032, d[01], c1132, quotient[22], s1131, c1131);
addsub a11_32(y[21], d[00], quotient[22], quotient[22], s1132, c1132);


addsub a12_00(s1101, d[32], c1201, quotient[21], s1200, quotient[20]);
addsub a12_01(s1102, d[31], c1202, quotient[21], s1201, c1201);
addsub a12_02(s1103, d[30], c1203, quotient[21], s1202, c1202);
addsub a12_03(s1104, d[29], c1204, quotient[21], s1203, c1203);
addsub a12_04(s1105, d[28], c1205, quotient[21], s1204, c1204);
addsub a12_05(s1106, d[27], c1206, quotient[21], s1205, c1205);
addsub a12_06(s1107, d[26], c1207, quotient[21], s1206, c1206);
addsub a12_07(s1108, d[25], c1208, quotient[21], s1207, c1207);
addsub a12_08(s1109, d[24], c1209, quotient[21], s1208, c1208);
addsub a12_09(s1110, d[23], c1210, quotient[21], s1209, c1209);
addsub a12_10(s1111, d[22], c1211, quotient[21], s1210, c1210);
addsub a12_11(s1112, d[21], c1212, quotient[21], s1211, c1211);
addsub a12_12(s1113, d[20], c1213, quotient[21], s1212, c1212);
addsub a12_13(s1114, d[19], c1214, quotient[21], s1213, c1213);
addsub a12_14(s1115, d[18], c1215, quotient[21], s1214, c1214);
addsub a12_15(s1116, d[17], c1216, quotient[21], s1215, c1215);
addsub a12_16(s1117, d[16], c1217, quotient[21], s1216, c1216);
addsub a12_17(s1118, d[15], c1218, quotient[21], s1217, c1217);
addsub a12_18(s1119, d[14], c1219, quotient[21], s1218, c1218);
addsub a12_19(s1120, d[13], c1220, quotient[21], s1219, c1219);
addsub a12_20(s1121, d[12], c1221, quotient[21], s1220, c1220);
addsub a12_21(s1122, d[11], c1222, quotient[21], s1221, c1221);
addsub a12_22(s1123, d[10], c1223, quotient[21], s1222, c1222);
addsub a12_23(s1124, d[09], c1224, quotient[21], s1223, c1223);
addsub a12_24(s1125, d[08], c1225, quotient[21], s1224, c1224);
addsub a12_25(s1126, d[07], c1226, quotient[21], s1225, c1225);
addsub a12_26(s1127, d[06], c1227, quotient[21], s1226, c1226);
addsub a12_27(s1128, d[05], c1228, quotient[21], s1227, c1227);
addsub a12_28(s1129, d[04], c1229, quotient[21], s1228, c1228);
addsub a12_29(s1130, d[03], c1230, quotient[21], s1229, c1229);
addsub a12_30(s1131, d[02], c1231, quotient[21], s1230, c1230);
addsub a12_31(s1132, d[01], c1232, quotient[21], s1231, c1231);
addsub a12_32(y[20], d[00], quotient[21], quotient[21], s1232, c1232);


addsub a13_00(s1201, d[32], c1301, quotient[20], s1300, quotient[19]);
addsub a13_01(s1202, d[31], c1302, quotient[20], s1301, c1301);
addsub a13_02(s1203, d[30], c1303, quotient[20], s1302, c1302);
addsub a13_03(s1204, d[29], c1304, quotient[20], s1303, c1303);
addsub a13_04(s1205, d[28], c1305, quotient[20], s1304, c1304);
addsub a13_05(s1206, d[27], c1306, quotient[20], s1305, c1305);
addsub a13_06(s1207, d[26], c1307, quotient[20], s1306, c1306);
addsub a13_07(s1208, d[25], c1308, quotient[20], s1307, c1307);
addsub a13_08(s1209, d[24], c1309, quotient[20], s1308, c1308);
addsub a13_09(s1210, d[23], c1310, quotient[20], s1309, c1309);
addsub a13_10(s1211, d[22], c1311, quotient[20], s1310, c1310);
addsub a13_11(s1212, d[21], c1312, quotient[20], s1311, c1311);
addsub a13_12(s1213, d[20], c1313, quotient[20], s1312, c1312);
addsub a13_13(s1214, d[19], c1314, quotient[20], s1313, c1313);
addsub a13_14(s1215, d[18], c1315, quotient[20], s1314, c1314);
addsub a13_15(s1216, d[17], c1316, quotient[20], s1315, c1315);
addsub a13_16(s1217, d[16], c1317, quotient[20], s1316, c1316);
addsub a13_17(s1218, d[15], c1318, quotient[20], s1317, c1317);
addsub a13_18(s1219, d[14], c1319, quotient[20], s1318, c1318);
addsub a13_19(s1220, d[13], c1320, quotient[20], s1319, c1319);
addsub a13_20(s1221, d[12], c1321, quotient[20], s1320, c1320);
addsub a13_21(s1222, d[11], c1322, quotient[20], s1321, c1321);
addsub a13_22(s1223, d[10], c1323, quotient[20], s1322, c1322);
addsub a13_23(s1224, d[09], c1324, quotient[20], s1323, c1323);
addsub a13_24(s1225, d[08], c1325, quotient[20], s1324, c1324);
addsub a13_25(s1226, d[07], c1326, quotient[20], s1325, c1325);
addsub a13_26(s1227, d[06], c1327, quotient[20], s1326, c1326);
addsub a13_27(s1228, d[05], c1328, quotient[20], s1327, c1327);
addsub a13_28(s1229, d[04], c1329, quotient[20], s1328, c1328);
addsub a13_29(s1230, d[03], c1330, quotient[20], s1329, c1329);
addsub a13_30(s1231, d[02], c1331, quotient[20], s1330, c1330);
addsub a13_31(s1232, d[01], c1332, quotient[20], s1331, c1331);
addsub a13_32(y[19], d[00], quotient[20], quotient[20], s1332, c1332);


addsub a14_00(s1301, d[32], c1401, quotient[19], s1400, quotient[18]);
addsub a14_01(s1302, d[31], c1402, quotient[19], s1401, c1401);
addsub a14_02(s1303, d[30], c1403, quotient[19], s1402, c1402);
addsub a14_03(s1304, d[29], c1404, quotient[19], s1403, c1403);
addsub a14_04(s1305, d[28], c1405, quotient[19], s1404, c1404);
addsub a14_05(s1306, d[27], c1406, quotient[19], s1405, c1405);
addsub a14_06(s1307, d[26], c1407, quotient[19], s1406, c1406);
addsub a14_07(s1308, d[25], c1408, quotient[19], s1407, c1407);
addsub a14_08(s1309, d[24], c1409, quotient[19], s1408, c1408);
addsub a14_09(s1310, d[23], c1410, quotient[19], s1409, c1409);
addsub a14_10(s1311, d[22], c1411, quotient[19], s1410, c1410);
addsub a14_11(s1312, d[21], c1412, quotient[19], s1411, c1411);
addsub a14_12(s1313, d[20], c1413, quotient[19], s1412, c1412);
addsub a14_13(s1314, d[19], c1414, quotient[19], s1413, c1413);
addsub a14_14(s1315, d[18], c1415, quotient[19], s1414, c1414);
addsub a14_15(s1316, d[17], c1416, quotient[19], s1415, c1415);
addsub a14_16(s1317, d[16], c1417, quotient[19], s1416, c1416);
addsub a14_17(s1318, d[15], c1418, quotient[19], s1417, c1417);
addsub a14_18(s1319, d[14], c1419, quotient[19], s1418, c1418);
addsub a14_19(s1320, d[13], c1420, quotient[19], s1419, c1419);
addsub a14_20(s1321, d[12], c1421, quotient[19], s1420, c1420);
addsub a14_21(s1322, d[11], c1422, quotient[19], s1421, c1421);
addsub a14_22(s1323, d[10], c1423, quotient[19], s1422, c1422);
addsub a14_23(s1324, d[09], c1424, quotient[19], s1423, c1423);
addsub a14_24(s1325, d[08], c1425, quotient[19], s1424, c1424);
addsub a14_25(s1326, d[07], c1426, quotient[19], s1425, c1425);
addsub a14_26(s1327, d[06], c1427, quotient[19], s1426, c1426);
addsub a14_27(s1328, d[05], c1428, quotient[19], s1427, c1427);
addsub a14_28(s1329, d[04], c1429, quotient[19], s1428, c1428);
addsub a14_29(s1330, d[03], c1430, quotient[19], s1429, c1429);
addsub a14_30(s1331, d[02], c1431, quotient[19], s1430, c1430);
addsub a14_31(s1332, d[01], c1432, quotient[19], s1431, c1431);
addsub a14_32(y[18], d[00], quotient[19], quotient[19], s1432, c1432);


addsub a15_00(s1401, d[32], c1501, quotient[18], s1500, quotient[17]);
addsub a15_01(s1402, d[31], c1502, quotient[18], s1501, c1501);
addsub a15_02(s1403, d[30], c1503, quotient[18], s1502, c1502);
addsub a15_03(s1404, d[29], c1504, quotient[18], s1503, c1503);
addsub a15_04(s1405, d[28], c1505, quotient[18], s1504, c1504);
addsub a15_05(s1406, d[27], c1506, quotient[18], s1505, c1505);
addsub a15_06(s1407, d[26], c1507, quotient[18], s1506, c1506);
addsub a15_07(s1408, d[25], c1508, quotient[18], s1507, c1507);
addsub a15_08(s1409, d[24], c1509, quotient[18], s1508, c1508);
addsub a15_09(s1410, d[23], c1510, quotient[18], s1509, c1509);
addsub a15_10(s1411, d[22], c1511, quotient[18], s1510, c1510);
addsub a15_11(s1412, d[21], c1512, quotient[18], s1511, c1511);
addsub a15_12(s1413, d[20], c1513, quotient[18], s1512, c1512);
addsub a15_13(s1414, d[19], c1514, quotient[18], s1513, c1513);
addsub a15_14(s1415, d[18], c1515, quotient[18], s1514, c1514);
addsub a15_15(s1416, d[17], c1516, quotient[18], s1515, c1515);
addsub a15_16(s1417, d[16], c1517, quotient[18], s1516, c1516);
addsub a15_17(s1418, d[15], c1518, quotient[18], s1517, c1517);
addsub a15_18(s1419, d[14], c1519, quotient[18], s1518, c1518);
addsub a15_19(s1420, d[13], c1520, quotient[18], s1519, c1519);
addsub a15_20(s1421, d[12], c1521, quotient[18], s1520, c1520);
addsub a15_21(s1422, d[11], c1522, quotient[18], s1521, c1521);
addsub a15_22(s1423, d[10], c1523, quotient[18], s1522, c1522);
addsub a15_23(s1424, d[09], c1524, quotient[18], s1523, c1523);
addsub a15_24(s1425, d[08], c1525, quotient[18], s1524, c1524);
addsub a15_25(s1426, d[07], c1526, quotient[18], s1525, c1525);
addsub a15_26(s1427, d[06], c1527, quotient[18], s1526, c1526);
addsub a15_27(s1428, d[05], c1528, quotient[18], s1527, c1527);
addsub a15_28(s1429, d[04], c1529, quotient[18], s1528, c1528);
addsub a15_29(s1430, d[03], c1530, quotient[18], s1529, c1529);
addsub a15_30(s1431, d[02], c1531, quotient[18], s1530, c1530);
addsub a15_31(s1432, d[01], c1532, quotient[18], s1531, c1531);
addsub a15_32(y[17], d[00], quotient[18], quotient[18], s1532, c1532);


addsub a16_00(s1501, d[32], c1601, quotient[17], s1600, quotient[16]);
addsub a16_01(s1502, d[31], c1602, quotient[17], s1601, c1601);
addsub a16_02(s1503, d[30], c1603, quotient[17], s1602, c1602);
addsub a16_03(s1504, d[29], c1604, quotient[17], s1603, c1603);
addsub a16_04(s1505, d[28], c1605, quotient[17], s1604, c1604);
addsub a16_05(s1506, d[27], c1606, quotient[17], s1605, c1605);
addsub a16_06(s1507, d[26], c1607, quotient[17], s1606, c1606);
addsub a16_07(s1508, d[25], c1608, quotient[17], s1607, c1607);
addsub a16_08(s1509, d[24], c1609, quotient[17], s1608, c1608);
addsub a16_09(s1510, d[23], c1610, quotient[17], s1609, c1609);
addsub a16_10(s1511, d[22], c1611, quotient[17], s1610, c1610);
addsub a16_11(s1512, d[21], c1612, quotient[17], s1611, c1611);
addsub a16_12(s1513, d[20], c1613, quotient[17], s1612, c1612);
addsub a16_13(s1514, d[19], c1614, quotient[17], s1613, c1613);
addsub a16_14(s1515, d[18], c1615, quotient[17], s1614, c1614);
addsub a16_15(s1516, d[17], c1616, quotient[17], s1615, c1615);
addsub a16_16(s1517, d[16], c1617, quotient[17], s1616, c1616);
addsub a16_17(s1518, d[15], c1618, quotient[17], s1617, c1617);
addsub a16_18(s1519, d[14], c1619, quotient[17], s1618, c1618);
addsub a16_19(s1520, d[13], c1620, quotient[17], s1619, c1619);
addsub a16_20(s1521, d[12], c1621, quotient[17], s1620, c1620);
addsub a16_21(s1522, d[11], c1622, quotient[17], s1621, c1621);
addsub a16_22(s1523, d[10], c1623, quotient[17], s1622, c1622);
addsub a16_23(s1524, d[09], c1624, quotient[17], s1623, c1623);
addsub a16_24(s1525, d[08], c1625, quotient[17], s1624, c1624);
addsub a16_25(s1526, d[07], c1626, quotient[17], s1625, c1625);
addsub a16_26(s1527, d[06], c1627, quotient[17], s1626, c1626);
addsub a16_27(s1528, d[05], c1628, quotient[17], s1627, c1627);
addsub a16_28(s1529, d[04], c1629, quotient[17], s1628, c1628);
addsub a16_29(s1530, d[03], c1630, quotient[17], s1629, c1629);
addsub a16_30(s1531, d[02], c1631, quotient[17], s1630, c1630);
addsub a16_31(s1532, d[01], c1632, quotient[17], s1631, c1631);
addsub a16_32(y[16], d[00], quotient[17], quotient[17], s1632, c1632);


addsub a17_00(s1601, d[32], c1701, quotient[16], s1700, quotient[15]);
addsub a17_01(s1602, d[31], c1702, quotient[16], s1701, c1701);
addsub a17_02(s1603, d[30], c1703, quotient[16], s1702, c1702);
addsub a17_03(s1604, d[29], c1704, quotient[16], s1703, c1703);
addsub a17_04(s1605, d[28], c1705, quotient[16], s1704, c1704);
addsub a17_05(s1606, d[27], c1706, quotient[16], s1705, c1705);
addsub a17_06(s1607, d[26], c1707, quotient[16], s1706, c1706);
addsub a17_07(s1608, d[25], c1708, quotient[16], s1707, c1707);
addsub a17_08(s1609, d[24], c1709, quotient[16], s1708, c1708);
addsub a17_09(s1610, d[23], c1710, quotient[16], s1709, c1709);
addsub a17_10(s1611, d[22], c1711, quotient[16], s1710, c1710);
addsub a17_11(s1612, d[21], c1712, quotient[16], s1711, c1711);
addsub a17_12(s1613, d[20], c1713, quotient[16], s1712, c1712);
addsub a17_13(s1614, d[19], c1714, quotient[16], s1713, c1713);
addsub a17_14(s1615, d[18], c1715, quotient[16], s1714, c1714);
addsub a17_15(s1616, d[17], c1716, quotient[16], s1715, c1715);
addsub a17_16(s1617, d[16], c1717, quotient[16], s1716, c1716);
addsub a17_17(s1618, d[15], c1718, quotient[16], s1717, c1717);
addsub a17_18(s1619, d[14], c1719, quotient[16], s1718, c1718);
addsub a17_19(s1620, d[13], c1720, quotient[16], s1719, c1719);
addsub a17_20(s1621, d[12], c1721, quotient[16], s1720, c1720);
addsub a17_21(s1622, d[11], c1722, quotient[16], s1721, c1721);
addsub a17_22(s1623, d[10], c1723, quotient[16], s1722, c1722);
addsub a17_23(s1624, d[09], c1724, quotient[16], s1723, c1723);
addsub a17_24(s1625, d[08], c1725, quotient[16], s1724, c1724);
addsub a17_25(s1626, d[07], c1726, quotient[16], s1725, c1725);
addsub a17_26(s1627, d[06], c1727, quotient[16], s1726, c1726);
addsub a17_27(s1628, d[05], c1728, quotient[16], s1727, c1727);
addsub a17_28(s1629, d[04], c1729, quotient[16], s1728, c1728);
addsub a17_29(s1630, d[03], c1730, quotient[16], s1729, c1729);
addsub a17_30(s1631, d[02], c1731, quotient[16], s1730, c1730);
addsub a17_31(s1632, d[01], c1732, quotient[16], s1731, c1731);
addsub a17_32(y[15], d[00], quotient[16], quotient[16], s1732, c1732);


addsub a18_00(s1701, d[32], c1801, quotient[15], s1800, quotient[14]);
addsub a18_01(s1702, d[31], c1802, quotient[15], s1801, c1801);
addsub a18_02(s1703, d[30], c1803, quotient[15], s1802, c1802);
addsub a18_03(s1704, d[29], c1804, quotient[15], s1803, c1803);
addsub a18_04(s1705, d[28], c1805, quotient[15], s1804, c1804);
addsub a18_05(s1706, d[27], c1806, quotient[15], s1805, c1805);
addsub a18_06(s1707, d[26], c1807, quotient[15], s1806, c1806);
addsub a18_07(s1708, d[25], c1808, quotient[15], s1807, c1807);
addsub a18_08(s1709, d[24], c1809, quotient[15], s1808, c1808);
addsub a18_09(s1710, d[23], c1810, quotient[15], s1809, c1809);
addsub a18_10(s1711, d[22], c1811, quotient[15], s1810, c1810);
addsub a18_11(s1712, d[21], c1812, quotient[15], s1811, c1811);
addsub a18_12(s1713, d[20], c1813, quotient[15], s1812, c1812);
addsub a18_13(s1714, d[19], c1814, quotient[15], s1813, c1813);
addsub a18_14(s1715, d[18], c1815, quotient[15], s1814, c1814);
addsub a18_15(s1716, d[17], c1816, quotient[15], s1815, c1815);
addsub a18_16(s1717, d[16], c1817, quotient[15], s1816, c1816);
addsub a18_17(s1718, d[15], c1818, quotient[15], s1817, c1817);
addsub a18_18(s1719, d[14], c1819, quotient[15], s1818, c1818);
addsub a18_19(s1720, d[13], c1820, quotient[15], s1819, c1819);
addsub a18_20(s1721, d[12], c1821, quotient[15], s1820, c1820);
addsub a18_21(s1722, d[11], c1822, quotient[15], s1821, c1821);
addsub a18_22(s1723, d[10], c1823, quotient[15], s1822, c1822);
addsub a18_23(s1724, d[09], c1824, quotient[15], s1823, c1823);
addsub a18_24(s1725, d[08], c1825, quotient[15], s1824, c1824);
addsub a18_25(s1726, d[07], c1826, quotient[15], s1825, c1825);
addsub a18_26(s1727, d[06], c1827, quotient[15], s1826, c1826);
addsub a18_27(s1728, d[05], c1828, quotient[15], s1827, c1827);
addsub a18_28(s1729, d[04], c1829, quotient[15], s1828, c1828);
addsub a18_29(s1730, d[03], c1830, quotient[15], s1829, c1829);
addsub a18_30(s1731, d[02], c1831, quotient[15], s1830, c1830);
addsub a18_31(s1732, d[01], c1832, quotient[15], s1831, c1831);
addsub a18_32(y[14], d[00], quotient[15], quotient[15], s1832, c1832);


addsub a19_00(s1801, d[32], c1901, quotient[14], s1900, quotient[13]);
addsub a19_01(s1802, d[31], c1902, quotient[14], s1901, c1901);
addsub a19_02(s1803, d[30], c1903, quotient[14], s1902, c1902);
addsub a19_03(s1804, d[29], c1904, quotient[14], s1903, c1903);
addsub a19_04(s1805, d[28], c1905, quotient[14], s1904, c1904);
addsub a19_05(s1806, d[27], c1906, quotient[14], s1905, c1905);
addsub a19_06(s1807, d[26], c1907, quotient[14], s1906, c1906);
addsub a19_07(s1808, d[25], c1908, quotient[14], s1907, c1907);
addsub a19_08(s1809, d[24], c1909, quotient[14], s1908, c1908);
addsub a19_09(s1810, d[23], c1910, quotient[14], s1909, c1909);
addsub a19_10(s1811, d[22], c1911, quotient[14], s1910, c1910);
addsub a19_11(s1812, d[21], c1912, quotient[14], s1911, c1911);
addsub a19_12(s1813, d[20], c1913, quotient[14], s1912, c1912);
addsub a19_13(s1814, d[19], c1914, quotient[14], s1913, c1913);
addsub a19_14(s1815, d[18], c1915, quotient[14], s1914, c1914);
addsub a19_15(s1816, d[17], c1916, quotient[14], s1915, c1915);
addsub a19_16(s1817, d[16], c1917, quotient[14], s1916, c1916);
addsub a19_17(s1818, d[15], c1918, quotient[14], s1917, c1917);
addsub a19_18(s1819, d[14], c1919, quotient[14], s1918, c1918);
addsub a19_19(s1820, d[13], c1920, quotient[14], s1919, c1919);
addsub a19_20(s1821, d[12], c1921, quotient[14], s1920, c1920);
addsub a19_21(s1822, d[11], c1922, quotient[14], s1921, c1921);
addsub a19_22(s1823, d[10], c1923, quotient[14], s1922, c1922);
addsub a19_23(s1824, d[09], c1924, quotient[14], s1923, c1923);
addsub a19_24(s1825, d[08], c1925, quotient[14], s1924, c1924);
addsub a19_25(s1826, d[07], c1926, quotient[14], s1925, c1925);
addsub a19_26(s1827, d[06], c1927, quotient[14], s1926, c1926);
addsub a19_27(s1828, d[05], c1928, quotient[14], s1927, c1927);
addsub a19_28(s1829, d[04], c1929, quotient[14], s1928, c1928);
addsub a19_29(s1830, d[03], c1930, quotient[14], s1929, c1929);
addsub a19_30(s1831, d[02], c1931, quotient[14], s1930, c1930);
addsub a19_31(s1832, d[01], c1932, quotient[14], s1931, c1931);
addsub a19_32(y[13], d[00], quotient[14], quotient[14], s1932, c1932);


addsub a20_00(s1901, d[32], c2001, quotient[13], s2000, quotient[12]);
addsub a20_01(s1902, d[31], c2002, quotient[13], s2001, c2001);
addsub a20_02(s1903, d[30], c2003, quotient[13], s2002, c2002);
addsub a20_03(s1904, d[29], c2004, quotient[13], s2003, c2003);
addsub a20_04(s1905, d[28], c2005, quotient[13], s2004, c2004);
addsub a20_05(s1906, d[27], c2006, quotient[13], s2005, c2005);
addsub a20_06(s1907, d[26], c2007, quotient[13], s2006, c2006);
addsub a20_07(s1908, d[25], c2008, quotient[13], s2007, c2007);
addsub a20_08(s1909, d[24], c2009, quotient[13], s2008, c2008);
addsub a20_09(s1910, d[23], c2010, quotient[13], s2009, c2009);
addsub a20_10(s1911, d[22], c2011, quotient[13], s2010, c2010);
addsub a20_11(s1912, d[21], c2012, quotient[13], s2011, c2011);
addsub a20_12(s1913, d[20], c2013, quotient[13], s2012, c2012);
addsub a20_13(s1914, d[19], c2014, quotient[13], s2013, c2013);
addsub a20_14(s1915, d[18], c2015, quotient[13], s2014, c2014);
addsub a20_15(s1916, d[17], c2016, quotient[13], s2015, c2015);
addsub a20_16(s1917, d[16], c2017, quotient[13], s2016, c2016);
addsub a20_17(s1918, d[15], c2018, quotient[13], s2017, c2017);
addsub a20_18(s1919, d[14], c2019, quotient[13], s2018, c2018);
addsub a20_19(s1920, d[13], c2020, quotient[13], s2019, c2019);
addsub a20_20(s1921, d[12], c2021, quotient[13], s2020, c2020);
addsub a20_21(s1922, d[11], c2022, quotient[13], s2021, c2021);
addsub a20_22(s1923, d[10], c2023, quotient[13], s2022, c2022);
addsub a20_23(s1924, d[09], c2024, quotient[13], s2023, c2023);
addsub a20_24(s1925, d[08], c2025, quotient[13], s2024, c2024);
addsub a20_25(s1926, d[07], c2026, quotient[13], s2025, c2025);
addsub a20_26(s1927, d[06], c2027, quotient[13], s2026, c2026);
addsub a20_27(s1928, d[05], c2028, quotient[13], s2027, c2027);
addsub a20_28(s1929, d[04], c2029, quotient[13], s2028, c2028);
addsub a20_29(s1930, d[03], c2030, quotient[13], s2029, c2029);
addsub a20_30(s1931, d[02], c2031, quotient[13], s2030, c2030);
addsub a20_31(s1932, d[01], c2032, quotient[13], s2031, c2031);
addsub a20_32(y[12], d[00], quotient[13], quotient[13], s2032, c2032);


addsub a21_00(s2001, d[32], c2101, quotient[12], s2100, quotient[11]);
addsub a21_01(s2002, d[31], c2102, quotient[12], s2101, c2101);
addsub a21_02(s2003, d[30], c2103, quotient[12], s2102, c2102);
addsub a21_03(s2004, d[29], c2104, quotient[12], s2103, c2103);
addsub a21_04(s2005, d[28], c2105, quotient[12], s2104, c2104);
addsub a21_05(s2006, d[27], c2106, quotient[12], s2105, c2105);
addsub a21_06(s2007, d[26], c2107, quotient[12], s2106, c2106);
addsub a21_07(s2008, d[25], c2108, quotient[12], s2107, c2107);
addsub a21_08(s2009, d[24], c2109, quotient[12], s2108, c2108);
addsub a21_09(s2010, d[23], c2110, quotient[12], s2109, c2109);
addsub a21_10(s2011, d[22], c2111, quotient[12], s2110, c2110);
addsub a21_11(s2012, d[21], c2112, quotient[12], s2111, c2111);
addsub a21_12(s2013, d[20], c2113, quotient[12], s2112, c2112);
addsub a21_13(s2014, d[19], c2114, quotient[12], s2113, c2113);
addsub a21_14(s2015, d[18], c2115, quotient[12], s2114, c2114);
addsub a21_15(s2016, d[17], c2116, quotient[12], s2115, c2115);
addsub a21_16(s2017, d[16], c2117, quotient[12], s2116, c2116);
addsub a21_17(s2018, d[15], c2118, quotient[12], s2117, c2117);
addsub a21_18(s2019, d[14], c2119, quotient[12], s2118, c2118);
addsub a21_19(s2020, d[13], c2120, quotient[12], s2119, c2119);
addsub a21_20(s2021, d[12], c2121, quotient[12], s2120, c2120);
addsub a21_21(s2022, d[11], c2122, quotient[12], s2121, c2121);
addsub a21_22(s2023, d[10], c2123, quotient[12], s2122, c2122);
addsub a21_23(s2024, d[09], c2124, quotient[12], s2123, c2123);
addsub a21_24(s2025, d[08], c2125, quotient[12], s2124, c2124);
addsub a21_25(s2026, d[07], c2126, quotient[12], s2125, c2125);
addsub a21_26(s2027, d[06], c2127, quotient[12], s2126, c2126);
addsub a21_27(s2028, d[05], c2128, quotient[12], s2127, c2127);
addsub a21_28(s2029, d[04], c2129, quotient[12], s2128, c2128);
addsub a21_29(s2030, d[03], c2130, quotient[12], s2129, c2129);
addsub a21_30(s2031, d[02], c2131, quotient[12], s2130, c2130);
addsub a21_31(s2032, d[01], c2132, quotient[12], s2131, c2131);
addsub a21_32(y[11], d[00], quotient[12], quotient[12], s2132, c2132);


addsub a22_00(s2101, d[32], c2201, quotient[11], s2200, quotient[10]);
addsub a22_01(s2102, d[31], c2202, quotient[11], s2201, c2201);
addsub a22_02(s2103, d[30], c2203, quotient[11], s2202, c2202);
addsub a22_03(s2104, d[29], c2204, quotient[11], s2203, c2203);
addsub a22_04(s2105, d[28], c2205, quotient[11], s2204, c2204);
addsub a22_05(s2106, d[27], c2206, quotient[11], s2205, c2205);
addsub a22_06(s2107, d[26], c2207, quotient[11], s2206, c2206);
addsub a22_07(s2108, d[25], c2208, quotient[11], s2207, c2207);
addsub a22_08(s2109, d[24], c2209, quotient[11], s2208, c2208);
addsub a22_09(s2110, d[23], c2210, quotient[11], s2209, c2209);
addsub a22_10(s2111, d[22], c2211, quotient[11], s2210, c2210);
addsub a22_11(s2112, d[21], c2212, quotient[11], s2211, c2211);
addsub a22_12(s2113, d[20], c2213, quotient[11], s2212, c2212);
addsub a22_13(s2114, d[19], c2214, quotient[11], s2213, c2213);
addsub a22_14(s2115, d[18], c2215, quotient[11], s2214, c2214);
addsub a22_15(s2116, d[17], c2216, quotient[11], s2215, c2215);
addsub a22_16(s2117, d[16], c2217, quotient[11], s2216, c2216);
addsub a22_17(s2118, d[15], c2218, quotient[11], s2217, c2217);
addsub a22_18(s2119, d[14], c2219, quotient[11], s2218, c2218);
addsub a22_19(s2120, d[13], c2220, quotient[11], s2219, c2219);
addsub a22_20(s2121, d[12], c2221, quotient[11], s2220, c2220);
addsub a22_21(s2122, d[11], c2222, quotient[11], s2221, c2221);
addsub a22_22(s2123, d[10], c2223, quotient[11], s2222, c2222);
addsub a22_23(s2124, d[09], c2224, quotient[11], s2223, c2223);
addsub a22_24(s2125, d[08], c2225, quotient[11], s2224, c2224);
addsub a22_25(s2126, d[07], c2226, quotient[11], s2225, c2225);
addsub a22_26(s2127, d[06], c2227, quotient[11], s2226, c2226);
addsub a22_27(s2128, d[05], c2228, quotient[11], s2227, c2227);
addsub a22_28(s2129, d[04], c2229, quotient[11], s2228, c2228);
addsub a22_29(s2130, d[03], c2230, quotient[11], s2229, c2229);
addsub a22_30(s2131, d[02], c2231, quotient[11], s2230, c2230);
addsub a22_31(s2132, d[01], c2232, quotient[11], s2231, c2231);
addsub a22_32(y[10], d[00], quotient[11], quotient[11], s2232, c2232);


addsub a23_00(s2201, d[32], c2301, quotient[10], s2300, quotient[09]);
addsub a23_01(s2202, d[31], c2302, quotient[10], s2301, c2301);
addsub a23_02(s2203, d[30], c2303, quotient[10], s2302, c2302);
addsub a23_03(s2204, d[29], c2304, quotient[10], s2303, c2303);
addsub a23_04(s2205, d[28], c2305, quotient[10], s2304, c2304);
addsub a23_05(s2206, d[27], c2306, quotient[10], s2305, c2305);
addsub a23_06(s2207, d[26], c2307, quotient[10], s2306, c2306);
addsub a23_07(s2208, d[25], c2308, quotient[10], s2307, c2307);
addsub a23_08(s2209, d[24], c2309, quotient[10], s2308, c2308);
addsub a23_09(s2210, d[23], c2310, quotient[10], s2309, c2309);
addsub a23_10(s2211, d[22], c2311, quotient[10], s2310, c2310);
addsub a23_11(s2212, d[21], c2312, quotient[10], s2311, c2311);
addsub a23_12(s2213, d[20], c2313, quotient[10], s2312, c2312);
addsub a23_13(s2214, d[19], c2314, quotient[10], s2313, c2313);
addsub a23_14(s2215, d[18], c2315, quotient[10], s2314, c2314);
addsub a23_15(s2216, d[17], c2316, quotient[10], s2315, c2315);
addsub a23_16(s2217, d[16], c2317, quotient[10], s2316, c2316);
addsub a23_17(s2218, d[15], c2318, quotient[10], s2317, c2317);
addsub a23_18(s2219, d[14], c2319, quotient[10], s2318, c2318);
addsub a23_19(s2220, d[13], c2320, quotient[10], s2319, c2319);
addsub a23_20(s2221, d[12], c2321, quotient[10], s2320, c2320);
addsub a23_21(s2222, d[11], c2322, quotient[10], s2321, c2321);
addsub a23_22(s2223, d[10], c2323, quotient[10], s2322, c2322);
addsub a23_23(s2224, d[09], c2324, quotient[10], s2323, c2323);
addsub a23_24(s2225, d[08], c2325, quotient[10], s2324, c2324);
addsub a23_25(s2226, d[07], c2326, quotient[10], s2325, c2325);
addsub a23_26(s2227, d[06], c2327, quotient[10], s2326, c2326);
addsub a23_27(s2228, d[05], c2328, quotient[10], s2327, c2327);
addsub a23_28(s2229, d[04], c2329, quotient[10], s2328, c2328);
addsub a23_29(s2230, d[03], c2330, quotient[10], s2329, c2329);
addsub a23_30(s2231, d[02], c2331, quotient[10], s2330, c2330);
addsub a23_31(s2232, d[01], c2332, quotient[10], s2331, c2331);
addsub a23_32(y[09], d[00], quotient[10], quotient[10], s2332, c2332);


addsub a24_00(s2301, d[32], c2401, quotient[09], s2400, quotient[08]);
addsub a24_01(s2302, d[31], c2402, quotient[09], s2401, c2401);
addsub a24_02(s2303, d[30], c2403, quotient[09], s2402, c2402);
addsub a24_03(s2304, d[29], c2404, quotient[09], s2403, c2403);
addsub a24_04(s2305, d[28], c2405, quotient[09], s2404, c2404);
addsub a24_05(s2306, d[27], c2406, quotient[09], s2405, c2405);
addsub a24_06(s2307, d[26], c2407, quotient[09], s2406, c2406);
addsub a24_07(s2308, d[25], c2408, quotient[09], s2407, c2407);
addsub a24_08(s2309, d[24], c2409, quotient[09], s2408, c2408);
addsub a24_09(s2310, d[23], c2410, quotient[09], s2409, c2409);
addsub a24_10(s2311, d[22], c2411, quotient[09], s2410, c2410);
addsub a24_11(s2312, d[21], c2412, quotient[09], s2411, c2411);
addsub a24_12(s2313, d[20], c2413, quotient[09], s2412, c2412);
addsub a24_13(s2314, d[19], c2414, quotient[09], s2413, c2413);
addsub a24_14(s2315, d[18], c2415, quotient[09], s2414, c2414);
addsub a24_15(s2316, d[17], c2416, quotient[09], s2415, c2415);
addsub a24_16(s2317, d[16], c2417, quotient[09], s2416, c2416);
addsub a24_17(s2318, d[15], c2418, quotient[09], s2417, c2417);
addsub a24_18(s2319, d[14], c2419, quotient[09], s2418, c2418);
addsub a24_19(s2320, d[13], c2420, quotient[09], s2419, c2419);
addsub a24_20(s2321, d[12], c2421, quotient[09], s2420, c2420);
addsub a24_21(s2322, d[11], c2422, quotient[09], s2421, c2421);
addsub a24_22(s2323, d[10], c2423, quotient[09], s2422, c2422);
addsub a24_23(s2324, d[09], c2424, quotient[09], s2423, c2423);
addsub a24_24(s2325, d[08], c2425, quotient[09], s2424, c2424);
addsub a24_25(s2326, d[07], c2426, quotient[09], s2425, c2425);
addsub a24_26(s2327, d[06], c2427, quotient[09], s2426, c2426);
addsub a24_27(s2328, d[05], c2428, quotient[09], s2427, c2427);
addsub a24_28(s2329, d[04], c2429, quotient[09], s2428, c2428);
addsub a24_29(s2330, d[03], c2430, quotient[09], s2429, c2429);
addsub a24_30(s2331, d[02], c2431, quotient[09], s2430, c2430);
addsub a24_31(s2332, d[01], c2432, quotient[09], s2431, c2431);
addsub a24_32(y[08], d[00], quotient[09], quotient[09], s2432, c2432);


addsub a25_00(s2401, d[32], c2501, quotient[08], s2500, quotient[07]);
addsub a25_01(s2402, d[31], c2502, quotient[08], s2501, c2501);
addsub a25_02(s2403, d[30], c2503, quotient[08], s2502, c2502);
addsub a25_03(s2404, d[29], c2504, quotient[08], s2503, c2503);
addsub a25_04(s2405, d[28], c2505, quotient[08], s2504, c2504);
addsub a25_05(s2406, d[27], c2506, quotient[08], s2505, c2505);
addsub a25_06(s2407, d[26], c2507, quotient[08], s2506, c2506);
addsub a25_07(s2408, d[25], c2508, quotient[08], s2507, c2507);
addsub a25_08(s2409, d[24], c2509, quotient[08], s2508, c2508);
addsub a25_09(s2410, d[23], c2510, quotient[08], s2509, c2509);
addsub a25_10(s2411, d[22], c2511, quotient[08], s2510, c2510);
addsub a25_11(s2412, d[21], c2512, quotient[08], s2511, c2511);
addsub a25_12(s2413, d[20], c2513, quotient[08], s2512, c2512);
addsub a25_13(s2414, d[19], c2514, quotient[08], s2513, c2513);
addsub a25_14(s2415, d[18], c2515, quotient[08], s2514, c2514);
addsub a25_15(s2416, d[17], c2516, quotient[08], s2515, c2515);
addsub a25_16(s2417, d[16], c2517, quotient[08], s2516, c2516);
addsub a25_17(s2418, d[15], c2518, quotient[08], s2517, c2517);
addsub a25_18(s2419, d[14], c2519, quotient[08], s2518, c2518);
addsub a25_19(s2420, d[13], c2520, quotient[08], s2519, c2519);
addsub a25_20(s2421, d[12], c2521, quotient[08], s2520, c2520);
addsub a25_21(s2422, d[11], c2522, quotient[08], s2521, c2521);
addsub a25_22(s2423, d[10], c2523, quotient[08], s2522, c2522);
addsub a25_23(s2424, d[09], c2524, quotient[08], s2523, c2523);
addsub a25_24(s2425, d[08], c2525, quotient[08], s2524, c2524);
addsub a25_25(s2426, d[07], c2526, quotient[08], s2525, c2525);
addsub a25_26(s2427, d[06], c2527, quotient[08], s2526, c2526);
addsub a25_27(s2428, d[05], c2528, quotient[08], s2527, c2527);
addsub a25_28(s2429, d[04], c2529, quotient[08], s2528, c2528);
addsub a25_29(s2430, d[03], c2530, quotient[08], s2529, c2529);
addsub a25_30(s2431, d[02], c2531, quotient[08], s2530, c2530);
addsub a25_31(s2432, d[01], c2532, quotient[08], s2531, c2531);
addsub a25_32(y[07], d[00], quotient[08], quotient[08], s2532, c2532);


addsub a26_00(s2501, d[32], c2601, quotient[07], s2600, quotient[06]);
addsub a26_01(s2502, d[31], c2602, quotient[07], s2601, c2601);
addsub a26_02(s2503, d[30], c2603, quotient[07], s2602, c2602);
addsub a26_03(s2504, d[29], c2604, quotient[07], s2603, c2603);
addsub a26_04(s2505, d[28], c2605, quotient[07], s2604, c2604);
addsub a26_05(s2506, d[27], c2606, quotient[07], s2605, c2605);
addsub a26_06(s2507, d[26], c2607, quotient[07], s2606, c2606);
addsub a26_07(s2508, d[25], c2608, quotient[07], s2607, c2607);
addsub a26_08(s2509, d[24], c2609, quotient[07], s2608, c2608);
addsub a26_09(s2510, d[23], c2610, quotient[07], s2609, c2609);
addsub a26_10(s2511, d[22], c2611, quotient[07], s2610, c2610);
addsub a26_11(s2512, d[21], c2612, quotient[07], s2611, c2611);
addsub a26_12(s2513, d[20], c2613, quotient[07], s2612, c2612);
addsub a26_13(s2514, d[19], c2614, quotient[07], s2613, c2613);
addsub a26_14(s2515, d[18], c2615, quotient[07], s2614, c2614);
addsub a26_15(s2516, d[17], c2616, quotient[07], s2615, c2615);
addsub a26_16(s2517, d[16], c2617, quotient[07], s2616, c2616);
addsub a26_17(s2518, d[15], c2618, quotient[07], s2617, c2617);
addsub a26_18(s2519, d[14], c2619, quotient[07], s2618, c2618);
addsub a26_19(s2520, d[13], c2620, quotient[07], s2619, c2619);
addsub a26_20(s2521, d[12], c2621, quotient[07], s2620, c2620);
addsub a26_21(s2522, d[11], c2622, quotient[07], s2621, c2621);
addsub a26_22(s2523, d[10], c2623, quotient[07], s2622, c2622);
addsub a26_23(s2524, d[09], c2624, quotient[07], s2623, c2623);
addsub a26_24(s2525, d[08], c2625, quotient[07], s2624, c2624);
addsub a26_25(s2526, d[07], c2626, quotient[07], s2625, c2625);
addsub a26_26(s2527, d[06], c2627, quotient[07], s2626, c2626);
addsub a26_27(s2528, d[05], c2628, quotient[07], s2627, c2627);
addsub a26_28(s2529, d[04], c2629, quotient[07], s2628, c2628);
addsub a26_29(s2530, d[03], c2630, quotient[07], s2629, c2629);
addsub a26_30(s2531, d[02], c2631, quotient[07], s2630, c2630);
addsub a26_31(s2532, d[01], c2632, quotient[07], s2631, c2631);
addsub a26_32(y[06], d[00], quotient[07], quotient[07], s2632, c2632);


addsub a27_00(s2601, d[32], c2701, quotient[06], s2700, quotient[05]);
addsub a27_01(s2602, d[31], c2702, quotient[06], s2701, c2701);
addsub a27_02(s2603, d[30], c2703, quotient[06], s2702, c2702);
addsub a27_03(s2604, d[29], c2704, quotient[06], s2703, c2703);
addsub a27_04(s2605, d[28], c2705, quotient[06], s2704, c2704);
addsub a27_05(s2606, d[27], c2706, quotient[06], s2705, c2705);
addsub a27_06(s2607, d[26], c2707, quotient[06], s2706, c2706);
addsub a27_07(s2608, d[25], c2708, quotient[06], s2707, c2707);
addsub a27_08(s2609, d[24], c2709, quotient[06], s2708, c2708);
addsub a27_09(s2610, d[23], c2710, quotient[06], s2709, c2709);
addsub a27_10(s2611, d[22], c2711, quotient[06], s2710, c2710);
addsub a27_11(s2612, d[21], c2712, quotient[06], s2711, c2711);
addsub a27_12(s2613, d[20], c2713, quotient[06], s2712, c2712);
addsub a27_13(s2614, d[19], c2714, quotient[06], s2713, c2713);
addsub a27_14(s2615, d[18], c2715, quotient[06], s2714, c2714);
addsub a27_15(s2616, d[17], c2716, quotient[06], s2715, c2715);
addsub a27_16(s2617, d[16], c2717, quotient[06], s2716, c2716);
addsub a27_17(s2618, d[15], c2718, quotient[06], s2717, c2717);
addsub a27_18(s2619, d[14], c2719, quotient[06], s2718, c2718);
addsub a27_19(s2620, d[13], c2720, quotient[06], s2719, c2719);
addsub a27_20(s2621, d[12], c2721, quotient[06], s2720, c2720);
addsub a27_21(s2622, d[11], c2722, quotient[06], s2721, c2721);
addsub a27_22(s2623, d[10], c2723, quotient[06], s2722, c2722);
addsub a27_23(s2624, d[09], c2724, quotient[06], s2723, c2723);
addsub a27_24(s2625, d[08], c2725, quotient[06], s2724, c2724);
addsub a27_25(s2626, d[07], c2726, quotient[06], s2725, c2725);
addsub a27_26(s2627, d[06], c2727, quotient[06], s2726, c2726);
addsub a27_27(s2628, d[05], c2728, quotient[06], s2727, c2727);
addsub a27_28(s2629, d[04], c2729, quotient[06], s2728, c2728);
addsub a27_29(s2630, d[03], c2730, quotient[06], s2729, c2729);
addsub a27_30(s2631, d[02], c2731, quotient[06], s2730, c2730);
addsub a27_31(s2632, d[01], c2732, quotient[06], s2731, c2731);
addsub a27_32(y[05], d[00], quotient[06], quotient[06], s2732, c2732);


addsub a28_00(s2701, d[32], c2801, quotient[05], s2800, quotient[04]);
addsub a28_01(s2702, d[31], c2802, quotient[05], s2801, c2801);
addsub a28_02(s2703, d[30], c2803, quotient[05], s2802, c2802);
addsub a28_03(s2704, d[29], c2804, quotient[05], s2803, c2803);
addsub a28_04(s2705, d[28], c2805, quotient[05], s2804, c2804);
addsub a28_05(s2706, d[27], c2806, quotient[05], s2805, c2805);
addsub a28_06(s2707, d[26], c2807, quotient[05], s2806, c2806);
addsub a28_07(s2708, d[25], c2808, quotient[05], s2807, c2807);
addsub a28_08(s2709, d[24], c2809, quotient[05], s2808, c2808);
addsub a28_09(s2710, d[23], c2810, quotient[05], s2809, c2809);
addsub a28_10(s2711, d[22], c2811, quotient[05], s2810, c2810);
addsub a28_11(s2712, d[21], c2812, quotient[05], s2811, c2811);
addsub a28_12(s2713, d[20], c2813, quotient[05], s2812, c2812);
addsub a28_13(s2714, d[19], c2814, quotient[05], s2813, c2813);
addsub a28_14(s2715, d[18], c2815, quotient[05], s2814, c2814);
addsub a28_15(s2716, d[17], c2816, quotient[05], s2815, c2815);
addsub a28_16(s2717, d[16], c2817, quotient[05], s2816, c2816);
addsub a28_17(s2718, d[15], c2818, quotient[05], s2817, c2817);
addsub a28_18(s2719, d[14], c2819, quotient[05], s2818, c2818);
addsub a28_19(s2720, d[13], c2820, quotient[05], s2819, c2819);
addsub a28_20(s2721, d[12], c2821, quotient[05], s2820, c2820);
addsub a28_21(s2722, d[11], c2822, quotient[05], s2821, c2821);
addsub a28_22(s2723, d[10], c2823, quotient[05], s2822, c2822);
addsub a28_23(s2724, d[09], c2824, quotient[05], s2823, c2823);
addsub a28_24(s2725, d[08], c2825, quotient[05], s2824, c2824);
addsub a28_25(s2726, d[07], c2826, quotient[05], s2825, c2825);
addsub a28_26(s2727, d[06], c2827, quotient[05], s2826, c2826);
addsub a28_27(s2728, d[05], c2828, quotient[05], s2827, c2827);
addsub a28_28(s2729, d[04], c2829, quotient[05], s2828, c2828);
addsub a28_29(s2730, d[03], c2830, quotient[05], s2829, c2829);
addsub a28_30(s2731, d[02], c2831, quotient[05], s2830, c2830);
addsub a28_31(s2732, d[01], c2832, quotient[05], s2831, c2831);
addsub a28_32(y[04], d[00], quotient[05], quotient[05], s2832, c2832);


addsub a29_00(s2801, d[32], c2901, quotient[04], s2900, quotient[03]);
addsub a29_01(s2802, d[31], c2902, quotient[04], s2901, c2901);
addsub a29_02(s2803, d[30], c2903, quotient[04], s2902, c2902);
addsub a29_03(s2804, d[29], c2904, quotient[04], s2903, c2903);
addsub a29_04(s2805, d[28], c2905, quotient[04], s2904, c2904);
addsub a29_05(s2806, d[27], c2906, quotient[04], s2905, c2905);
addsub a29_06(s2807, d[26], c2907, quotient[04], s2906, c2906);
addsub a29_07(s2808, d[25], c2908, quotient[04], s2907, c2907);
addsub a29_08(s2809, d[24], c2909, quotient[04], s2908, c2908);
addsub a29_09(s2810, d[23], c2910, quotient[04], s2909, c2909);
addsub a29_10(s2811, d[22], c2911, quotient[04], s2910, c2910);
addsub a29_11(s2812, d[21], c2912, quotient[04], s2911, c2911);
addsub a29_12(s2813, d[20], c2913, quotient[04], s2912, c2912);
addsub a29_13(s2814, d[19], c2914, quotient[04], s2913, c2913);
addsub a29_14(s2815, d[18], c2915, quotient[04], s2914, c2914);
addsub a29_15(s2816, d[17], c2916, quotient[04], s2915, c2915);
addsub a29_16(s2817, d[16], c2917, quotient[04], s2916, c2916);
addsub a29_17(s2818, d[15], c2918, quotient[04], s2917, c2917);
addsub a29_18(s2819, d[14], c2919, quotient[04], s2918, c2918);
addsub a29_19(s2820, d[13], c2920, quotient[04], s2919, c2919);
addsub a29_20(s2821, d[12], c2921, quotient[04], s2920, c2920);
addsub a29_21(s2822, d[11], c2922, quotient[04], s2921, c2921);
addsub a29_22(s2823, d[10], c2923, quotient[04], s2922, c2922);
addsub a29_23(s2824, d[09], c2924, quotient[04], s2923, c2923);
addsub a29_24(s2825, d[08], c2925, quotient[04], s2924, c2924);
addsub a29_25(s2826, d[07], c2926, quotient[04], s2925, c2925);
addsub a29_26(s2827, d[06], c2927, quotient[04], s2926, c2926);
addsub a29_27(s2828, d[05], c2928, quotient[04], s2927, c2927);
addsub a29_28(s2829, d[04], c2929, quotient[04], s2928, c2928);
addsub a29_29(s2830, d[03], c2930, quotient[04], s2929, c2929);
addsub a29_30(s2831, d[02], c2931, quotient[04], s2930, c2930);
addsub a29_31(s2832, d[01], c2932, quotient[04], s2931, c2931);
addsub a29_32(y[03], d[00], quotient[04], quotient[04], s2932, c2932);


addsub a30_00(s2901, d[32], c3001, quotient[03], s3000, quotient[02]);
addsub a30_01(s2902, d[31], c3002, quotient[03], s3001, c3001);
addsub a30_02(s2903, d[30], c3003, quotient[03], s3002, c3002);
addsub a30_03(s2904, d[29], c3004, quotient[03], s3003, c3003);
addsub a30_04(s2905, d[28], c3005, quotient[03], s3004, c3004);
addsub a30_05(s2906, d[27], c3006, quotient[03], s3005, c3005);
addsub a30_06(s2907, d[26], c3007, quotient[03], s3006, c3006);
addsub a30_07(s2908, d[25], c3008, quotient[03], s3007, c3007);
addsub a30_08(s2909, d[24], c3009, quotient[03], s3008, c3008);
addsub a30_09(s2910, d[23], c3010, quotient[03], s3009, c3009);
addsub a30_10(s2911, d[22], c3011, quotient[03], s3010, c3010);
addsub a30_11(s2912, d[21], c3012, quotient[03], s3011, c3011);
addsub a30_12(s2913, d[20], c3013, quotient[03], s3012, c3012);
addsub a30_13(s2914, d[19], c3014, quotient[03], s3013, c3013);
addsub a30_14(s2915, d[18], c3015, quotient[03], s3014, c3014);
addsub a30_15(s2916, d[17], c3016, quotient[03], s3015, c3015);
addsub a30_16(s2917, d[16], c3017, quotient[03], s3016, c3016);
addsub a30_17(s2918, d[15], c3018, quotient[03], s3017, c3017);
addsub a30_18(s2919, d[14], c3019, quotient[03], s3018, c3018);
addsub a30_19(s2920, d[13], c3020, quotient[03], s3019, c3019);
addsub a30_20(s2921, d[12], c3021, quotient[03], s3020, c3020);
addsub a30_21(s2922, d[11], c3022, quotient[03], s3021, c3021);
addsub a30_22(s2923, d[10], c3023, quotient[03], s3022, c3022);
addsub a30_23(s2924, d[09], c3024, quotient[03], s3023, c3023);
addsub a30_24(s2925, d[08], c3025, quotient[03], s3024, c3024);
addsub a30_25(s2926, d[07], c3026, quotient[03], s3025, c3025);
addsub a30_26(s2927, d[06], c3027, quotient[03], s3026, c3026);
addsub a30_27(s2928, d[05], c3028, quotient[03], s3027, c3027);
addsub a30_28(s2929, d[04], c3029, quotient[03], s3028, c3028);
addsub a30_29(s2930, d[03], c3030, quotient[03], s3029, c3029);
addsub a30_30(s2931, d[02], c3031, quotient[03], s3030, c3030);
addsub a30_31(s2932, d[01], c3032, quotient[03], s3031, c3031);
addsub a30_32(y[02], d[00], quotient[03], quotient[03], s3032, c3032);


addsub a31_00(s3001, d[32], c3101, quotient[02], s3100, quotient[01]);
addsub a31_01(s3002, d[31], c3102, quotient[02], s3101, c3101);
addsub a31_02(s3003, d[30], c3103, quotient[02], s3102, c3102);
addsub a31_03(s3004, d[29], c3104, quotient[02], s3103, c3103);
addsub a31_04(s3005, d[28], c3105, quotient[02], s3104, c3104);
addsub a31_05(s3006, d[27], c3106, quotient[02], s3105, c3105);
addsub a31_06(s3007, d[26], c3107, quotient[02], s3106, c3106);
addsub a31_07(s3008, d[25], c3108, quotient[02], s3107, c3107);
addsub a31_08(s3009, d[24], c3109, quotient[02], s3108, c3108);
addsub a31_09(s3010, d[23], c3110, quotient[02], s3109, c3109);
addsub a31_10(s3011, d[22], c3111, quotient[02], s3110, c3110);
addsub a31_11(s3012, d[21], c3112, quotient[02], s3111, c3111);
addsub a31_12(s3013, d[20], c3113, quotient[02], s3112, c3112);
addsub a31_13(s3014, d[19], c3114, quotient[02], s3113, c3113);
addsub a31_14(s3015, d[18], c3115, quotient[02], s3114, c3114);
addsub a31_15(s3016, d[17], c3116, quotient[02], s3115, c3115);
addsub a31_16(s3017, d[16], c3117, quotient[02], s3116, c3116);
addsub a31_17(s3018, d[15], c3118, quotient[02], s3117, c3117);
addsub a31_18(s3019, d[14], c3119, quotient[02], s3118, c3118);
addsub a31_19(s3020, d[13], c3120, quotient[02], s3119, c3119);
addsub a31_20(s3021, d[12], c3121, quotient[02], s3120, c3120);
addsub a31_21(s3022, d[11], c3122, quotient[02], s3121, c3121);
addsub a31_22(s3023, d[10], c3123, quotient[02], s3122, c3122);
addsub a31_23(s3024, d[09], c3124, quotient[02], s3123, c3123);
addsub a31_24(s3025, d[08], c3125, quotient[02], s3124, c3124);
addsub a31_25(s3026, d[07], c3126, quotient[02], s3125, c3125);
addsub a31_26(s3027, d[06], c3127, quotient[02], s3126, c3126);
addsub a31_27(s3028, d[05], c3128, quotient[02], s3127, c3127);
addsub a31_28(s3029, d[04], c3129, quotient[02], s3128, c3128);
addsub a31_29(s3030, d[03], c3130, quotient[02], s3129, c3129);
addsub a31_30(s3031, d[02], c3131, quotient[02], s3130, c3130);
addsub a31_31(s3032, d[01], c3132, quotient[02], s3131, c3131);
addsub a31_32(y[01], d[00], quotient[02], quotient[02], s3132, c3132);


addsub a32_00(s3101, d[32], c3201, quotient[01], s3200, quotient[00]);
addsub a32_01(s3102, d[31], c3202, quotient[01], s3201, c3201);
addsub a32_02(s3103, d[30], c3203, quotient[01], s3202, c3202);
addsub a32_03(s3104, d[29], c3204, quotient[01], s3203, c3203);
addsub a32_04(s3105, d[28], c3205, quotient[01], s3204, c3204);
addsub a32_05(s3106, d[27], c3206, quotient[01], s3205, c3205);
addsub a32_06(s3107, d[26], c3207, quotient[01], s3206, c3206);
addsub a32_07(s3108, d[25], c3208, quotient[01], s3207, c3207);
addsub a32_08(s3109, d[24], c3209, quotient[01], s3208, c3208);
addsub a32_09(s3110, d[23], c3210, quotient[01], s3209, c3209);
addsub a32_10(s3111, d[22], c3211, quotient[01], s3210, c3210);
addsub a32_11(s3112, d[21], c3212, quotient[01], s3211, c3211);
addsub a32_12(s3113, d[20], c3213, quotient[01], s3212, c3212);
addsub a32_13(s3114, d[19], c3214, quotient[01], s3213, c3213);
addsub a32_14(s3115, d[18], c3215, quotient[01], s3214, c3214);
addsub a32_15(s3116, d[17], c3216, quotient[01], s3215, c3215);
addsub a32_16(s3117, d[16], c3217, quotient[01], s3216, c3216);
addsub a32_17(s3118, d[15], c3218, quotient[01], s3217, c3217);
addsub a32_18(s3119, d[14], c3219, quotient[01], s3218, c3218);
addsub a32_19(s3120, d[13], c3220, quotient[01], s3219, c3219);
addsub a32_20(s3121, d[12], c3221, quotient[01], s3220, c3220);
addsub a32_21(s3122, d[11], c3222, quotient[01], s3221, c3221);
addsub a32_22(s3123, d[10], c3223, quotient[01], s3222, c3222);
addsub a32_23(s3124, d[09], c3224, quotient[01], s3223, c3223);
addsub a32_24(s3125, d[08], c3225, quotient[01], s3224, c3224);
addsub a32_25(s3126, d[07], c3226, quotient[01], s3225, c3225);
addsub a32_26(s3127, d[06], c3227, quotient[01], s3226, c3226);
addsub a32_27(s3128, d[05], c3228, quotient[01], s3227, c3227);
addsub a32_28(s3129, d[04], c3229, quotient[01], s3228, c3228);
addsub a32_29(s3130, d[03], c3230, quotient[01], s3229, c3229);
addsub a32_30(s3131, d[02], c3231, quotient[01], s3230, c3230);
addsub a32_31(s3132, d[01], c3232, quotient[01], s3231, c3231);
addsub a32_32(y[00], d[00], quotient[01], quotient[01], s3232, c3232);


assign remainder = s3200 ? {s3200,s3201,s3202,s3203,s3204,s3205,s3206,s3207,s3208,s3209,s3210,s3211,s3212,s3213,s3214,s3215,s3216,s3217,s3218,s3219,s3220,s3221,s3222,s3223,s3224,s3225,s3226,s3227,s3228,s3229,s3230,s3231,s3232} + divisor : {s3200,s3201,s3202,s3203,s3204,s3205,s3206,s3207,s3208,s3209,s3210,s3211,s3212,s3213,s3214,s3215,s3216,s3217,s3218,s3219,s3220,s3221,s3222,s3223,s3224,s3225,s3226,s3227,s3228,s3229,s3230,s3231,s3232};

always @(posedge clk) begin
    if (rst) begin
        y <= { 32'b0, dividend };
        d <= { 1'b0, divisor };
    end
end
endmodule
