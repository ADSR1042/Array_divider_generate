module divider_24bit(
    input wire clk,
    input wire rst,
    input wire [23:0] dividend,
    input wire [23:0] divisor,
    output wire [24:0] quotient,
    output wire [24:0] remainder
);
wire c0001,c0002,c0003,c0004,c0005,c0006,c0007,c0008,c0009,c0010,c0011,c0012,c0013,c0014,c0015,c0016,c0017,c0018,c0019,c0020,c0021,c0022,c0023,c0024;
wire c0101,c0102,c0103,c0104,c0105,c0106,c0107,c0108,c0109,c0110,c0111,c0112,c0113,c0114,c0115,c0116,c0117,c0118,c0119,c0120,c0121,c0122,c0123,c0124;
wire c0201,c0202,c0203,c0204,c0205,c0206,c0207,c0208,c0209,c0210,c0211,c0212,c0213,c0214,c0215,c0216,c0217,c0218,c0219,c0220,c0221,c0222,c0223,c0224;
wire c0301,c0302,c0303,c0304,c0305,c0306,c0307,c0308,c0309,c0310,c0311,c0312,c0313,c0314,c0315,c0316,c0317,c0318,c0319,c0320,c0321,c0322,c0323,c0324;
wire c0401,c0402,c0403,c0404,c0405,c0406,c0407,c0408,c0409,c0410,c0411,c0412,c0413,c0414,c0415,c0416,c0417,c0418,c0419,c0420,c0421,c0422,c0423,c0424;
wire c0501,c0502,c0503,c0504,c0505,c0506,c0507,c0508,c0509,c0510,c0511,c0512,c0513,c0514,c0515,c0516,c0517,c0518,c0519,c0520,c0521,c0522,c0523,c0524;
wire c0601,c0602,c0603,c0604,c0605,c0606,c0607,c0608,c0609,c0610,c0611,c0612,c0613,c0614,c0615,c0616,c0617,c0618,c0619,c0620,c0621,c0622,c0623,c0624;
wire c0701,c0702,c0703,c0704,c0705,c0706,c0707,c0708,c0709,c0710,c0711,c0712,c0713,c0714,c0715,c0716,c0717,c0718,c0719,c0720,c0721,c0722,c0723,c0724;
wire c0801,c0802,c0803,c0804,c0805,c0806,c0807,c0808,c0809,c0810,c0811,c0812,c0813,c0814,c0815,c0816,c0817,c0818,c0819,c0820,c0821,c0822,c0823,c0824;
wire c0901,c0902,c0903,c0904,c0905,c0906,c0907,c0908,c0909,c0910,c0911,c0912,c0913,c0914,c0915,c0916,c0917,c0918,c0919,c0920,c0921,c0922,c0923,c0924;
wire c1001,c1002,c1003,c1004,c1005,c1006,c1007,c1008,c1009,c1010,c1011,c1012,c1013,c1014,c1015,c1016,c1017,c1018,c1019,c1020,c1021,c1022,c1023,c1024;
wire c1101,c1102,c1103,c1104,c1105,c1106,c1107,c1108,c1109,c1110,c1111,c1112,c1113,c1114,c1115,c1116,c1117,c1118,c1119,c1120,c1121,c1122,c1123,c1124;
wire c1201,c1202,c1203,c1204,c1205,c1206,c1207,c1208,c1209,c1210,c1211,c1212,c1213,c1214,c1215,c1216,c1217,c1218,c1219,c1220,c1221,c1222,c1223,c1224;
wire c1301,c1302,c1303,c1304,c1305,c1306,c1307,c1308,c1309,c1310,c1311,c1312,c1313,c1314,c1315,c1316,c1317,c1318,c1319,c1320,c1321,c1322,c1323,c1324;
wire c1401,c1402,c1403,c1404,c1405,c1406,c1407,c1408,c1409,c1410,c1411,c1412,c1413,c1414,c1415,c1416,c1417,c1418,c1419,c1420,c1421,c1422,c1423,c1424;
wire c1501,c1502,c1503,c1504,c1505,c1506,c1507,c1508,c1509,c1510,c1511,c1512,c1513,c1514,c1515,c1516,c1517,c1518,c1519,c1520,c1521,c1522,c1523,c1524;
wire c1601,c1602,c1603,c1604,c1605,c1606,c1607,c1608,c1609,c1610,c1611,c1612,c1613,c1614,c1615,c1616,c1617,c1618,c1619,c1620,c1621,c1622,c1623,c1624;
wire c1701,c1702,c1703,c1704,c1705,c1706,c1707,c1708,c1709,c1710,c1711,c1712,c1713,c1714,c1715,c1716,c1717,c1718,c1719,c1720,c1721,c1722,c1723,c1724;
wire c1801,c1802,c1803,c1804,c1805,c1806,c1807,c1808,c1809,c1810,c1811,c1812,c1813,c1814,c1815,c1816,c1817,c1818,c1819,c1820,c1821,c1822,c1823,c1824;
wire c1901,c1902,c1903,c1904,c1905,c1906,c1907,c1908,c1909,c1910,c1911,c1912,c1913,c1914,c1915,c1916,c1917,c1918,c1919,c1920,c1921,c1922,c1923,c1924;
wire c2001,c2002,c2003,c2004,c2005,c2006,c2007,c2008,c2009,c2010,c2011,c2012,c2013,c2014,c2015,c2016,c2017,c2018,c2019,c2020,c2021,c2022,c2023,c2024;
wire c2101,c2102,c2103,c2104,c2105,c2106,c2107,c2108,c2109,c2110,c2111,c2112,c2113,c2114,c2115,c2116,c2117,c2118,c2119,c2120,c2121,c2122,c2123,c2124;
wire c2201,c2202,c2203,c2204,c2205,c2206,c2207,c2208,c2209,c2210,c2211,c2212,c2213,c2214,c2215,c2216,c2217,c2218,c2219,c2220,c2221,c2222,c2223,c2224;
wire c2301,c2302,c2303,c2304,c2305,c2306,c2307,c2308,c2309,c2310,c2311,c2312,c2313,c2314,c2315,c2316,c2317,c2318,c2319,c2320,c2321,c2322,c2323,c2324;
wire c2401,c2402,c2403,c2404,c2405,c2406,c2407,c2408,c2409,c2410,c2411,c2412,c2413,c2414,c2415,c2416,c2417,c2418,c2419,c2420,c2421,c2422,c2423,c2424;
wire s0000,s0001,s0002,s0003,s0004,s0005,s0006,s0007,s0008,s0009,s0010,s0011,s0012,s0013,s0014,s0015,s0016,s0017,s0018,s0019,s0020,s0021,s0022,s0023,s0024;
wire s0100,s0101,s0102,s0103,s0104,s0105,s0106,s0107,s0108,s0109,s0110,s0111,s0112,s0113,s0114,s0115,s0116,s0117,s0118,s0119,s0120,s0121,s0122,s0123,s0124;
wire s0200,s0201,s0202,s0203,s0204,s0205,s0206,s0207,s0208,s0209,s0210,s0211,s0212,s0213,s0214,s0215,s0216,s0217,s0218,s0219,s0220,s0221,s0222,s0223,s0224;
wire s0300,s0301,s0302,s0303,s0304,s0305,s0306,s0307,s0308,s0309,s0310,s0311,s0312,s0313,s0314,s0315,s0316,s0317,s0318,s0319,s0320,s0321,s0322,s0323,s0324;
wire s0400,s0401,s0402,s0403,s0404,s0405,s0406,s0407,s0408,s0409,s0410,s0411,s0412,s0413,s0414,s0415,s0416,s0417,s0418,s0419,s0420,s0421,s0422,s0423,s0424;
wire s0500,s0501,s0502,s0503,s0504,s0505,s0506,s0507,s0508,s0509,s0510,s0511,s0512,s0513,s0514,s0515,s0516,s0517,s0518,s0519,s0520,s0521,s0522,s0523,s0524;
wire s0600,s0601,s0602,s0603,s0604,s0605,s0606,s0607,s0608,s0609,s0610,s0611,s0612,s0613,s0614,s0615,s0616,s0617,s0618,s0619,s0620,s0621,s0622,s0623,s0624;
wire s0700,s0701,s0702,s0703,s0704,s0705,s0706,s0707,s0708,s0709,s0710,s0711,s0712,s0713,s0714,s0715,s0716,s0717,s0718,s0719,s0720,s0721,s0722,s0723,s0724;
wire s0800,s0801,s0802,s0803,s0804,s0805,s0806,s0807,s0808,s0809,s0810,s0811,s0812,s0813,s0814,s0815,s0816,s0817,s0818,s0819,s0820,s0821,s0822,s0823,s0824;
wire s0900,s0901,s0902,s0903,s0904,s0905,s0906,s0907,s0908,s0909,s0910,s0911,s0912,s0913,s0914,s0915,s0916,s0917,s0918,s0919,s0920,s0921,s0922,s0923,s0924;
wire s1000,s1001,s1002,s1003,s1004,s1005,s1006,s1007,s1008,s1009,s1010,s1011,s1012,s1013,s1014,s1015,s1016,s1017,s1018,s1019,s1020,s1021,s1022,s1023,s1024;
wire s1100,s1101,s1102,s1103,s1104,s1105,s1106,s1107,s1108,s1109,s1110,s1111,s1112,s1113,s1114,s1115,s1116,s1117,s1118,s1119,s1120,s1121,s1122,s1123,s1124;
wire s1200,s1201,s1202,s1203,s1204,s1205,s1206,s1207,s1208,s1209,s1210,s1211,s1212,s1213,s1214,s1215,s1216,s1217,s1218,s1219,s1220,s1221,s1222,s1223,s1224;
wire s1300,s1301,s1302,s1303,s1304,s1305,s1306,s1307,s1308,s1309,s1310,s1311,s1312,s1313,s1314,s1315,s1316,s1317,s1318,s1319,s1320,s1321,s1322,s1323,s1324;
wire s1400,s1401,s1402,s1403,s1404,s1405,s1406,s1407,s1408,s1409,s1410,s1411,s1412,s1413,s1414,s1415,s1416,s1417,s1418,s1419,s1420,s1421,s1422,s1423,s1424;
wire s1500,s1501,s1502,s1503,s1504,s1505,s1506,s1507,s1508,s1509,s1510,s1511,s1512,s1513,s1514,s1515,s1516,s1517,s1518,s1519,s1520,s1521,s1522,s1523,s1524;
wire s1600,s1601,s1602,s1603,s1604,s1605,s1606,s1607,s1608,s1609,s1610,s1611,s1612,s1613,s1614,s1615,s1616,s1617,s1618,s1619,s1620,s1621,s1622,s1623,s1624;
wire s1700,s1701,s1702,s1703,s1704,s1705,s1706,s1707,s1708,s1709,s1710,s1711,s1712,s1713,s1714,s1715,s1716,s1717,s1718,s1719,s1720,s1721,s1722,s1723,s1724;
wire s1800,s1801,s1802,s1803,s1804,s1805,s1806,s1807,s1808,s1809,s1810,s1811,s1812,s1813,s1814,s1815,s1816,s1817,s1818,s1819,s1820,s1821,s1822,s1823,s1824;
wire s1900,s1901,s1902,s1903,s1904,s1905,s1906,s1907,s1908,s1909,s1910,s1911,s1912,s1913,s1914,s1915,s1916,s1917,s1918,s1919,s1920,s1921,s1922,s1923,s1924;
wire s2000,s2001,s2002,s2003,s2004,s2005,s2006,s2007,s2008,s2009,s2010,s2011,s2012,s2013,s2014,s2015,s2016,s2017,s2018,s2019,s2020,s2021,s2022,s2023,s2024;
wire s2100,s2101,s2102,s2103,s2104,s2105,s2106,s2107,s2108,s2109,s2110,s2111,s2112,s2113,s2114,s2115,s2116,s2117,s2118,s2119,s2120,s2121,s2122,s2123,s2124;
wire s2200,s2201,s2202,s2203,s2204,s2205,s2206,s2207,s2208,s2209,s2210,s2211,s2212,s2213,s2214,s2215,s2216,s2217,s2218,s2219,s2220,s2221,s2222,s2223,s2224;
wire s2300,s2301,s2302,s2303,s2304,s2305,s2306,s2307,s2308,s2309,s2310,s2311,s2312,s2313,s2314,s2315,s2316,s2317,s2318,s2319,s2320,s2321,s2322,s2323,s2324;
wire s2400,s2401,s2402,s2403,s2404,s2405,s2406,s2407,s2408,s2409,s2410,s2411,s2412,s2413,s2414,s2415,s2416,s2417,s2418,s2419,s2420,s2421,s2422,s2423,s2424;

reg [48:0] y;
reg [24:0] d;

addsub a0_00(y[48], d[24], c0001, 1'b1, s0000, quotient[24]);
addsub a0_01(y[47], d[23], c0002, 1'b1, s0001, c0001);
addsub a0_02(y[46], d[22], c0003, 1'b1, s0002, c0002);
addsub a0_03(y[45], d[21], c0004, 1'b1, s0003, c0003);
addsub a0_04(y[44], d[20], c0005, 1'b1, s0004, c0004);
addsub a0_05(y[43], d[19], c0006, 1'b1, s0005, c0005);
addsub a0_06(y[42], d[18], c0007, 1'b1, s0006, c0006);
addsub a0_07(y[41], d[17], c0008, 1'b1, s0007, c0007);
addsub a0_08(y[40], d[16], c0009, 1'b1, s0008, c0008);
addsub a0_09(y[39], d[15], c0010, 1'b1, s0009, c0009);
addsub a0_10(y[38], d[14], c0011, 1'b1, s0010, c0010);
addsub a0_11(y[37], d[13], c0012, 1'b1, s0011, c0011);
addsub a0_12(y[36], d[12], c0013, 1'b1, s0012, c0012);
addsub a0_13(y[35], d[11], c0014, 1'b1, s0013, c0013);
addsub a0_14(y[34], d[10], c0015, 1'b1, s0014, c0014);
addsub a0_15(y[33], d[09], c0016, 1'b1, s0015, c0015);
addsub a0_16(y[32], d[08], c0017, 1'b1, s0016, c0016);
addsub a0_17(y[31], d[07], c0018, 1'b1, s0017, c0017);
addsub a0_18(y[30], d[06], c0019, 1'b1, s0018, c0018);
addsub a0_19(y[29], d[05], c0020, 1'b1, s0019, c0019);
addsub a0_20(y[28], d[04], c0021, 1'b1, s0020, c0020);
addsub a0_21(y[27], d[03], c0022, 1'b1, s0021, c0021);
addsub a0_22(y[26], d[02], c0023, 1'b1, s0022, c0022);
addsub a0_23(y[25], d[01], c0024, 1'b1, s0023, c0023);
addsub a0_24(y[24], d[00], 1'b1, 1'b1, s0024, c0024);


addsub a01_00(s0001, d[24], c0101, quotient[24], s0100, quotient[23]);
addsub a01_01(s0002, d[23], c0102, quotient[24], s0101, c0101);
addsub a01_02(s0003, d[22], c0103, quotient[24], s0102, c0102);
addsub a01_03(s0004, d[21], c0104, quotient[24], s0103, c0103);
addsub a01_04(s0005, d[20], c0105, quotient[24], s0104, c0104);
addsub a01_05(s0006, d[19], c0106, quotient[24], s0105, c0105);
addsub a01_06(s0007, d[18], c0107, quotient[24], s0106, c0106);
addsub a01_07(s0008, d[17], c0108, quotient[24], s0107, c0107);
addsub a01_08(s0009, d[16], c0109, quotient[24], s0108, c0108);
addsub a01_09(s0010, d[15], c0110, quotient[24], s0109, c0109);
addsub a01_10(s0011, d[14], c0111, quotient[24], s0110, c0110);
addsub a01_11(s0012, d[13], c0112, quotient[24], s0111, c0111);
addsub a01_12(s0013, d[12], c0113, quotient[24], s0112, c0112);
addsub a01_13(s0014, d[11], c0114, quotient[24], s0113, c0113);
addsub a01_14(s0015, d[10], c0115, quotient[24], s0114, c0114);
addsub a01_15(s0016, d[09], c0116, quotient[24], s0115, c0115);
addsub a01_16(s0017, d[08], c0117, quotient[24], s0116, c0116);
addsub a01_17(s0018, d[07], c0118, quotient[24], s0117, c0117);
addsub a01_18(s0019, d[06], c0119, quotient[24], s0118, c0118);
addsub a01_19(s0020, d[05], c0120, quotient[24], s0119, c0119);
addsub a01_20(s0021, d[04], c0121, quotient[24], s0120, c0120);
addsub a01_21(s0022, d[03], c0122, quotient[24], s0121, c0121);
addsub a01_22(s0023, d[02], c0123, quotient[24], s0122, c0122);
addsub a01_23(s0024, d[01], c0124, quotient[24], s0123, c0123);
addsub a01_24(y[23], d[00], quotient[24], quotient[24], s0124, c0124);


addsub a02_00(s0101, d[24], c0201, quotient[23], s0200, quotient[22]);
addsub a02_01(s0102, d[23], c0202, quotient[23], s0201, c0201);
addsub a02_02(s0103, d[22], c0203, quotient[23], s0202, c0202);
addsub a02_03(s0104, d[21], c0204, quotient[23], s0203, c0203);
addsub a02_04(s0105, d[20], c0205, quotient[23], s0204, c0204);
addsub a02_05(s0106, d[19], c0206, quotient[23], s0205, c0205);
addsub a02_06(s0107, d[18], c0207, quotient[23], s0206, c0206);
addsub a02_07(s0108, d[17], c0208, quotient[23], s0207, c0207);
addsub a02_08(s0109, d[16], c0209, quotient[23], s0208, c0208);
addsub a02_09(s0110, d[15], c0210, quotient[23], s0209, c0209);
addsub a02_10(s0111, d[14], c0211, quotient[23], s0210, c0210);
addsub a02_11(s0112, d[13], c0212, quotient[23], s0211, c0211);
addsub a02_12(s0113, d[12], c0213, quotient[23], s0212, c0212);
addsub a02_13(s0114, d[11], c0214, quotient[23], s0213, c0213);
addsub a02_14(s0115, d[10], c0215, quotient[23], s0214, c0214);
addsub a02_15(s0116, d[09], c0216, quotient[23], s0215, c0215);
addsub a02_16(s0117, d[08], c0217, quotient[23], s0216, c0216);
addsub a02_17(s0118, d[07], c0218, quotient[23], s0217, c0217);
addsub a02_18(s0119, d[06], c0219, quotient[23], s0218, c0218);
addsub a02_19(s0120, d[05], c0220, quotient[23], s0219, c0219);
addsub a02_20(s0121, d[04], c0221, quotient[23], s0220, c0220);
addsub a02_21(s0122, d[03], c0222, quotient[23], s0221, c0221);
addsub a02_22(s0123, d[02], c0223, quotient[23], s0222, c0222);
addsub a02_23(s0124, d[01], c0224, quotient[23], s0223, c0223);
addsub a02_24(y[22], d[00], quotient[23], quotient[23], s0224, c0224);


addsub a03_00(s0201, d[24], c0301, quotient[22], s0300, quotient[21]);
addsub a03_01(s0202, d[23], c0302, quotient[22], s0301, c0301);
addsub a03_02(s0203, d[22], c0303, quotient[22], s0302, c0302);
addsub a03_03(s0204, d[21], c0304, quotient[22], s0303, c0303);
addsub a03_04(s0205, d[20], c0305, quotient[22], s0304, c0304);
addsub a03_05(s0206, d[19], c0306, quotient[22], s0305, c0305);
addsub a03_06(s0207, d[18], c0307, quotient[22], s0306, c0306);
addsub a03_07(s0208, d[17], c0308, quotient[22], s0307, c0307);
addsub a03_08(s0209, d[16], c0309, quotient[22], s0308, c0308);
addsub a03_09(s0210, d[15], c0310, quotient[22], s0309, c0309);
addsub a03_10(s0211, d[14], c0311, quotient[22], s0310, c0310);
addsub a03_11(s0212, d[13], c0312, quotient[22], s0311, c0311);
addsub a03_12(s0213, d[12], c0313, quotient[22], s0312, c0312);
addsub a03_13(s0214, d[11], c0314, quotient[22], s0313, c0313);
addsub a03_14(s0215, d[10], c0315, quotient[22], s0314, c0314);
addsub a03_15(s0216, d[09], c0316, quotient[22], s0315, c0315);
addsub a03_16(s0217, d[08], c0317, quotient[22], s0316, c0316);
addsub a03_17(s0218, d[07], c0318, quotient[22], s0317, c0317);
addsub a03_18(s0219, d[06], c0319, quotient[22], s0318, c0318);
addsub a03_19(s0220, d[05], c0320, quotient[22], s0319, c0319);
addsub a03_20(s0221, d[04], c0321, quotient[22], s0320, c0320);
addsub a03_21(s0222, d[03], c0322, quotient[22], s0321, c0321);
addsub a03_22(s0223, d[02], c0323, quotient[22], s0322, c0322);
addsub a03_23(s0224, d[01], c0324, quotient[22], s0323, c0323);
addsub a03_24(y[21], d[00], quotient[22], quotient[22], s0324, c0324);


addsub a04_00(s0301, d[24], c0401, quotient[21], s0400, quotient[20]);
addsub a04_01(s0302, d[23], c0402, quotient[21], s0401, c0401);
addsub a04_02(s0303, d[22], c0403, quotient[21], s0402, c0402);
addsub a04_03(s0304, d[21], c0404, quotient[21], s0403, c0403);
addsub a04_04(s0305, d[20], c0405, quotient[21], s0404, c0404);
addsub a04_05(s0306, d[19], c0406, quotient[21], s0405, c0405);
addsub a04_06(s0307, d[18], c0407, quotient[21], s0406, c0406);
addsub a04_07(s0308, d[17], c0408, quotient[21], s0407, c0407);
addsub a04_08(s0309, d[16], c0409, quotient[21], s0408, c0408);
addsub a04_09(s0310, d[15], c0410, quotient[21], s0409, c0409);
addsub a04_10(s0311, d[14], c0411, quotient[21], s0410, c0410);
addsub a04_11(s0312, d[13], c0412, quotient[21], s0411, c0411);
addsub a04_12(s0313, d[12], c0413, quotient[21], s0412, c0412);
addsub a04_13(s0314, d[11], c0414, quotient[21], s0413, c0413);
addsub a04_14(s0315, d[10], c0415, quotient[21], s0414, c0414);
addsub a04_15(s0316, d[09], c0416, quotient[21], s0415, c0415);
addsub a04_16(s0317, d[08], c0417, quotient[21], s0416, c0416);
addsub a04_17(s0318, d[07], c0418, quotient[21], s0417, c0417);
addsub a04_18(s0319, d[06], c0419, quotient[21], s0418, c0418);
addsub a04_19(s0320, d[05], c0420, quotient[21], s0419, c0419);
addsub a04_20(s0321, d[04], c0421, quotient[21], s0420, c0420);
addsub a04_21(s0322, d[03], c0422, quotient[21], s0421, c0421);
addsub a04_22(s0323, d[02], c0423, quotient[21], s0422, c0422);
addsub a04_23(s0324, d[01], c0424, quotient[21], s0423, c0423);
addsub a04_24(y[20], d[00], quotient[21], quotient[21], s0424, c0424);


addsub a05_00(s0401, d[24], c0501, quotient[20], s0500, quotient[19]);
addsub a05_01(s0402, d[23], c0502, quotient[20], s0501, c0501);
addsub a05_02(s0403, d[22], c0503, quotient[20], s0502, c0502);
addsub a05_03(s0404, d[21], c0504, quotient[20], s0503, c0503);
addsub a05_04(s0405, d[20], c0505, quotient[20], s0504, c0504);
addsub a05_05(s0406, d[19], c0506, quotient[20], s0505, c0505);
addsub a05_06(s0407, d[18], c0507, quotient[20], s0506, c0506);
addsub a05_07(s0408, d[17], c0508, quotient[20], s0507, c0507);
addsub a05_08(s0409, d[16], c0509, quotient[20], s0508, c0508);
addsub a05_09(s0410, d[15], c0510, quotient[20], s0509, c0509);
addsub a05_10(s0411, d[14], c0511, quotient[20], s0510, c0510);
addsub a05_11(s0412, d[13], c0512, quotient[20], s0511, c0511);
addsub a05_12(s0413, d[12], c0513, quotient[20], s0512, c0512);
addsub a05_13(s0414, d[11], c0514, quotient[20], s0513, c0513);
addsub a05_14(s0415, d[10], c0515, quotient[20], s0514, c0514);
addsub a05_15(s0416, d[09], c0516, quotient[20], s0515, c0515);
addsub a05_16(s0417, d[08], c0517, quotient[20], s0516, c0516);
addsub a05_17(s0418, d[07], c0518, quotient[20], s0517, c0517);
addsub a05_18(s0419, d[06], c0519, quotient[20], s0518, c0518);
addsub a05_19(s0420, d[05], c0520, quotient[20], s0519, c0519);
addsub a05_20(s0421, d[04], c0521, quotient[20], s0520, c0520);
addsub a05_21(s0422, d[03], c0522, quotient[20], s0521, c0521);
addsub a05_22(s0423, d[02], c0523, quotient[20], s0522, c0522);
addsub a05_23(s0424, d[01], c0524, quotient[20], s0523, c0523);
addsub a05_24(y[19], d[00], quotient[20], quotient[20], s0524, c0524);


addsub a06_00(s0501, d[24], c0601, quotient[19], s0600, quotient[18]);
addsub a06_01(s0502, d[23], c0602, quotient[19], s0601, c0601);
addsub a06_02(s0503, d[22], c0603, quotient[19], s0602, c0602);
addsub a06_03(s0504, d[21], c0604, quotient[19], s0603, c0603);
addsub a06_04(s0505, d[20], c0605, quotient[19], s0604, c0604);
addsub a06_05(s0506, d[19], c0606, quotient[19], s0605, c0605);
addsub a06_06(s0507, d[18], c0607, quotient[19], s0606, c0606);
addsub a06_07(s0508, d[17], c0608, quotient[19], s0607, c0607);
addsub a06_08(s0509, d[16], c0609, quotient[19], s0608, c0608);
addsub a06_09(s0510, d[15], c0610, quotient[19], s0609, c0609);
addsub a06_10(s0511, d[14], c0611, quotient[19], s0610, c0610);
addsub a06_11(s0512, d[13], c0612, quotient[19], s0611, c0611);
addsub a06_12(s0513, d[12], c0613, quotient[19], s0612, c0612);
addsub a06_13(s0514, d[11], c0614, quotient[19], s0613, c0613);
addsub a06_14(s0515, d[10], c0615, quotient[19], s0614, c0614);
addsub a06_15(s0516, d[09], c0616, quotient[19], s0615, c0615);
addsub a06_16(s0517, d[08], c0617, quotient[19], s0616, c0616);
addsub a06_17(s0518, d[07], c0618, quotient[19], s0617, c0617);
addsub a06_18(s0519, d[06], c0619, quotient[19], s0618, c0618);
addsub a06_19(s0520, d[05], c0620, quotient[19], s0619, c0619);
addsub a06_20(s0521, d[04], c0621, quotient[19], s0620, c0620);
addsub a06_21(s0522, d[03], c0622, quotient[19], s0621, c0621);
addsub a06_22(s0523, d[02], c0623, quotient[19], s0622, c0622);
addsub a06_23(s0524, d[01], c0624, quotient[19], s0623, c0623);
addsub a06_24(y[18], d[00], quotient[19], quotient[19], s0624, c0624);


addsub a07_00(s0601, d[24], c0701, quotient[18], s0700, quotient[17]);
addsub a07_01(s0602, d[23], c0702, quotient[18], s0701, c0701);
addsub a07_02(s0603, d[22], c0703, quotient[18], s0702, c0702);
addsub a07_03(s0604, d[21], c0704, quotient[18], s0703, c0703);
addsub a07_04(s0605, d[20], c0705, quotient[18], s0704, c0704);
addsub a07_05(s0606, d[19], c0706, quotient[18], s0705, c0705);
addsub a07_06(s0607, d[18], c0707, quotient[18], s0706, c0706);
addsub a07_07(s0608, d[17], c0708, quotient[18], s0707, c0707);
addsub a07_08(s0609, d[16], c0709, quotient[18], s0708, c0708);
addsub a07_09(s0610, d[15], c0710, quotient[18], s0709, c0709);
addsub a07_10(s0611, d[14], c0711, quotient[18], s0710, c0710);
addsub a07_11(s0612, d[13], c0712, quotient[18], s0711, c0711);
addsub a07_12(s0613, d[12], c0713, quotient[18], s0712, c0712);
addsub a07_13(s0614, d[11], c0714, quotient[18], s0713, c0713);
addsub a07_14(s0615, d[10], c0715, quotient[18], s0714, c0714);
addsub a07_15(s0616, d[09], c0716, quotient[18], s0715, c0715);
addsub a07_16(s0617, d[08], c0717, quotient[18], s0716, c0716);
addsub a07_17(s0618, d[07], c0718, quotient[18], s0717, c0717);
addsub a07_18(s0619, d[06], c0719, quotient[18], s0718, c0718);
addsub a07_19(s0620, d[05], c0720, quotient[18], s0719, c0719);
addsub a07_20(s0621, d[04], c0721, quotient[18], s0720, c0720);
addsub a07_21(s0622, d[03], c0722, quotient[18], s0721, c0721);
addsub a07_22(s0623, d[02], c0723, quotient[18], s0722, c0722);
addsub a07_23(s0624, d[01], c0724, quotient[18], s0723, c0723);
addsub a07_24(y[17], d[00], quotient[18], quotient[18], s0724, c0724);


addsub a08_00(s0701, d[24], c0801, quotient[17], s0800, quotient[16]);
addsub a08_01(s0702, d[23], c0802, quotient[17], s0801, c0801);
addsub a08_02(s0703, d[22], c0803, quotient[17], s0802, c0802);
addsub a08_03(s0704, d[21], c0804, quotient[17], s0803, c0803);
addsub a08_04(s0705, d[20], c0805, quotient[17], s0804, c0804);
addsub a08_05(s0706, d[19], c0806, quotient[17], s0805, c0805);
addsub a08_06(s0707, d[18], c0807, quotient[17], s0806, c0806);
addsub a08_07(s0708, d[17], c0808, quotient[17], s0807, c0807);
addsub a08_08(s0709, d[16], c0809, quotient[17], s0808, c0808);
addsub a08_09(s0710, d[15], c0810, quotient[17], s0809, c0809);
addsub a08_10(s0711, d[14], c0811, quotient[17], s0810, c0810);
addsub a08_11(s0712, d[13], c0812, quotient[17], s0811, c0811);
addsub a08_12(s0713, d[12], c0813, quotient[17], s0812, c0812);
addsub a08_13(s0714, d[11], c0814, quotient[17], s0813, c0813);
addsub a08_14(s0715, d[10], c0815, quotient[17], s0814, c0814);
addsub a08_15(s0716, d[09], c0816, quotient[17], s0815, c0815);
addsub a08_16(s0717, d[08], c0817, quotient[17], s0816, c0816);
addsub a08_17(s0718, d[07], c0818, quotient[17], s0817, c0817);
addsub a08_18(s0719, d[06], c0819, quotient[17], s0818, c0818);
addsub a08_19(s0720, d[05], c0820, quotient[17], s0819, c0819);
addsub a08_20(s0721, d[04], c0821, quotient[17], s0820, c0820);
addsub a08_21(s0722, d[03], c0822, quotient[17], s0821, c0821);
addsub a08_22(s0723, d[02], c0823, quotient[17], s0822, c0822);
addsub a08_23(s0724, d[01], c0824, quotient[17], s0823, c0823);
addsub a08_24(y[16], d[00], quotient[17], quotient[17], s0824, c0824);


addsub a09_00(s0801, d[24], c0901, quotient[16], s0900, quotient[15]);
addsub a09_01(s0802, d[23], c0902, quotient[16], s0901, c0901);
addsub a09_02(s0803, d[22], c0903, quotient[16], s0902, c0902);
addsub a09_03(s0804, d[21], c0904, quotient[16], s0903, c0903);
addsub a09_04(s0805, d[20], c0905, quotient[16], s0904, c0904);
addsub a09_05(s0806, d[19], c0906, quotient[16], s0905, c0905);
addsub a09_06(s0807, d[18], c0907, quotient[16], s0906, c0906);
addsub a09_07(s0808, d[17], c0908, quotient[16], s0907, c0907);
addsub a09_08(s0809, d[16], c0909, quotient[16], s0908, c0908);
addsub a09_09(s0810, d[15], c0910, quotient[16], s0909, c0909);
addsub a09_10(s0811, d[14], c0911, quotient[16], s0910, c0910);
addsub a09_11(s0812, d[13], c0912, quotient[16], s0911, c0911);
addsub a09_12(s0813, d[12], c0913, quotient[16], s0912, c0912);
addsub a09_13(s0814, d[11], c0914, quotient[16], s0913, c0913);
addsub a09_14(s0815, d[10], c0915, quotient[16], s0914, c0914);
addsub a09_15(s0816, d[09], c0916, quotient[16], s0915, c0915);
addsub a09_16(s0817, d[08], c0917, quotient[16], s0916, c0916);
addsub a09_17(s0818, d[07], c0918, quotient[16], s0917, c0917);
addsub a09_18(s0819, d[06], c0919, quotient[16], s0918, c0918);
addsub a09_19(s0820, d[05], c0920, quotient[16], s0919, c0919);
addsub a09_20(s0821, d[04], c0921, quotient[16], s0920, c0920);
addsub a09_21(s0822, d[03], c0922, quotient[16], s0921, c0921);
addsub a09_22(s0823, d[02], c0923, quotient[16], s0922, c0922);
addsub a09_23(s0824, d[01], c0924, quotient[16], s0923, c0923);
addsub a09_24(y[15], d[00], quotient[16], quotient[16], s0924, c0924);


addsub a10_00(s0901, d[24], c1001, quotient[15], s1000, quotient[14]);
addsub a10_01(s0902, d[23], c1002, quotient[15], s1001, c1001);
addsub a10_02(s0903, d[22], c1003, quotient[15], s1002, c1002);
addsub a10_03(s0904, d[21], c1004, quotient[15], s1003, c1003);
addsub a10_04(s0905, d[20], c1005, quotient[15], s1004, c1004);
addsub a10_05(s0906, d[19], c1006, quotient[15], s1005, c1005);
addsub a10_06(s0907, d[18], c1007, quotient[15], s1006, c1006);
addsub a10_07(s0908, d[17], c1008, quotient[15], s1007, c1007);
addsub a10_08(s0909, d[16], c1009, quotient[15], s1008, c1008);
addsub a10_09(s0910, d[15], c1010, quotient[15], s1009, c1009);
addsub a10_10(s0911, d[14], c1011, quotient[15], s1010, c1010);
addsub a10_11(s0912, d[13], c1012, quotient[15], s1011, c1011);
addsub a10_12(s0913, d[12], c1013, quotient[15], s1012, c1012);
addsub a10_13(s0914, d[11], c1014, quotient[15], s1013, c1013);
addsub a10_14(s0915, d[10], c1015, quotient[15], s1014, c1014);
addsub a10_15(s0916, d[09], c1016, quotient[15], s1015, c1015);
addsub a10_16(s0917, d[08], c1017, quotient[15], s1016, c1016);
addsub a10_17(s0918, d[07], c1018, quotient[15], s1017, c1017);
addsub a10_18(s0919, d[06], c1019, quotient[15], s1018, c1018);
addsub a10_19(s0920, d[05], c1020, quotient[15], s1019, c1019);
addsub a10_20(s0921, d[04], c1021, quotient[15], s1020, c1020);
addsub a10_21(s0922, d[03], c1022, quotient[15], s1021, c1021);
addsub a10_22(s0923, d[02], c1023, quotient[15], s1022, c1022);
addsub a10_23(s0924, d[01], c1024, quotient[15], s1023, c1023);
addsub a10_24(y[14], d[00], quotient[15], quotient[15], s1024, c1024);


addsub a11_00(s1001, d[24], c1101, quotient[14], s1100, quotient[13]);
addsub a11_01(s1002, d[23], c1102, quotient[14], s1101, c1101);
addsub a11_02(s1003, d[22], c1103, quotient[14], s1102, c1102);
addsub a11_03(s1004, d[21], c1104, quotient[14], s1103, c1103);
addsub a11_04(s1005, d[20], c1105, quotient[14], s1104, c1104);
addsub a11_05(s1006, d[19], c1106, quotient[14], s1105, c1105);
addsub a11_06(s1007, d[18], c1107, quotient[14], s1106, c1106);
addsub a11_07(s1008, d[17], c1108, quotient[14], s1107, c1107);
addsub a11_08(s1009, d[16], c1109, quotient[14], s1108, c1108);
addsub a11_09(s1010, d[15], c1110, quotient[14], s1109, c1109);
addsub a11_10(s1011, d[14], c1111, quotient[14], s1110, c1110);
addsub a11_11(s1012, d[13], c1112, quotient[14], s1111, c1111);
addsub a11_12(s1013, d[12], c1113, quotient[14], s1112, c1112);
addsub a11_13(s1014, d[11], c1114, quotient[14], s1113, c1113);
addsub a11_14(s1015, d[10], c1115, quotient[14], s1114, c1114);
addsub a11_15(s1016, d[09], c1116, quotient[14], s1115, c1115);
addsub a11_16(s1017, d[08], c1117, quotient[14], s1116, c1116);
addsub a11_17(s1018, d[07], c1118, quotient[14], s1117, c1117);
addsub a11_18(s1019, d[06], c1119, quotient[14], s1118, c1118);
addsub a11_19(s1020, d[05], c1120, quotient[14], s1119, c1119);
addsub a11_20(s1021, d[04], c1121, quotient[14], s1120, c1120);
addsub a11_21(s1022, d[03], c1122, quotient[14], s1121, c1121);
addsub a11_22(s1023, d[02], c1123, quotient[14], s1122, c1122);
addsub a11_23(s1024, d[01], c1124, quotient[14], s1123, c1123);
addsub a11_24(y[13], d[00], quotient[14], quotient[14], s1124, c1124);


addsub a12_00(s1101, d[24], c1201, quotient[13], s1200, quotient[12]);
addsub a12_01(s1102, d[23], c1202, quotient[13], s1201, c1201);
addsub a12_02(s1103, d[22], c1203, quotient[13], s1202, c1202);
addsub a12_03(s1104, d[21], c1204, quotient[13], s1203, c1203);
addsub a12_04(s1105, d[20], c1205, quotient[13], s1204, c1204);
addsub a12_05(s1106, d[19], c1206, quotient[13], s1205, c1205);
addsub a12_06(s1107, d[18], c1207, quotient[13], s1206, c1206);
addsub a12_07(s1108, d[17], c1208, quotient[13], s1207, c1207);
addsub a12_08(s1109, d[16], c1209, quotient[13], s1208, c1208);
addsub a12_09(s1110, d[15], c1210, quotient[13], s1209, c1209);
addsub a12_10(s1111, d[14], c1211, quotient[13], s1210, c1210);
addsub a12_11(s1112, d[13], c1212, quotient[13], s1211, c1211);
addsub a12_12(s1113, d[12], c1213, quotient[13], s1212, c1212);
addsub a12_13(s1114, d[11], c1214, quotient[13], s1213, c1213);
addsub a12_14(s1115, d[10], c1215, quotient[13], s1214, c1214);
addsub a12_15(s1116, d[09], c1216, quotient[13], s1215, c1215);
addsub a12_16(s1117, d[08], c1217, quotient[13], s1216, c1216);
addsub a12_17(s1118, d[07], c1218, quotient[13], s1217, c1217);
addsub a12_18(s1119, d[06], c1219, quotient[13], s1218, c1218);
addsub a12_19(s1120, d[05], c1220, quotient[13], s1219, c1219);
addsub a12_20(s1121, d[04], c1221, quotient[13], s1220, c1220);
addsub a12_21(s1122, d[03], c1222, quotient[13], s1221, c1221);
addsub a12_22(s1123, d[02], c1223, quotient[13], s1222, c1222);
addsub a12_23(s1124, d[01], c1224, quotient[13], s1223, c1223);
addsub a12_24(y[12], d[00], quotient[13], quotient[13], s1224, c1224);


addsub a13_00(s1201, d[24], c1301, quotient[12], s1300, quotient[11]);
addsub a13_01(s1202, d[23], c1302, quotient[12], s1301, c1301);
addsub a13_02(s1203, d[22], c1303, quotient[12], s1302, c1302);
addsub a13_03(s1204, d[21], c1304, quotient[12], s1303, c1303);
addsub a13_04(s1205, d[20], c1305, quotient[12], s1304, c1304);
addsub a13_05(s1206, d[19], c1306, quotient[12], s1305, c1305);
addsub a13_06(s1207, d[18], c1307, quotient[12], s1306, c1306);
addsub a13_07(s1208, d[17], c1308, quotient[12], s1307, c1307);
addsub a13_08(s1209, d[16], c1309, quotient[12], s1308, c1308);
addsub a13_09(s1210, d[15], c1310, quotient[12], s1309, c1309);
addsub a13_10(s1211, d[14], c1311, quotient[12], s1310, c1310);
addsub a13_11(s1212, d[13], c1312, quotient[12], s1311, c1311);
addsub a13_12(s1213, d[12], c1313, quotient[12], s1312, c1312);
addsub a13_13(s1214, d[11], c1314, quotient[12], s1313, c1313);
addsub a13_14(s1215, d[10], c1315, quotient[12], s1314, c1314);
addsub a13_15(s1216, d[09], c1316, quotient[12], s1315, c1315);
addsub a13_16(s1217, d[08], c1317, quotient[12], s1316, c1316);
addsub a13_17(s1218, d[07], c1318, quotient[12], s1317, c1317);
addsub a13_18(s1219, d[06], c1319, quotient[12], s1318, c1318);
addsub a13_19(s1220, d[05], c1320, quotient[12], s1319, c1319);
addsub a13_20(s1221, d[04], c1321, quotient[12], s1320, c1320);
addsub a13_21(s1222, d[03], c1322, quotient[12], s1321, c1321);
addsub a13_22(s1223, d[02], c1323, quotient[12], s1322, c1322);
addsub a13_23(s1224, d[01], c1324, quotient[12], s1323, c1323);
addsub a13_24(y[11], d[00], quotient[12], quotient[12], s1324, c1324);


addsub a14_00(s1301, d[24], c1401, quotient[11], s1400, quotient[10]);
addsub a14_01(s1302, d[23], c1402, quotient[11], s1401, c1401);
addsub a14_02(s1303, d[22], c1403, quotient[11], s1402, c1402);
addsub a14_03(s1304, d[21], c1404, quotient[11], s1403, c1403);
addsub a14_04(s1305, d[20], c1405, quotient[11], s1404, c1404);
addsub a14_05(s1306, d[19], c1406, quotient[11], s1405, c1405);
addsub a14_06(s1307, d[18], c1407, quotient[11], s1406, c1406);
addsub a14_07(s1308, d[17], c1408, quotient[11], s1407, c1407);
addsub a14_08(s1309, d[16], c1409, quotient[11], s1408, c1408);
addsub a14_09(s1310, d[15], c1410, quotient[11], s1409, c1409);
addsub a14_10(s1311, d[14], c1411, quotient[11], s1410, c1410);
addsub a14_11(s1312, d[13], c1412, quotient[11], s1411, c1411);
addsub a14_12(s1313, d[12], c1413, quotient[11], s1412, c1412);
addsub a14_13(s1314, d[11], c1414, quotient[11], s1413, c1413);
addsub a14_14(s1315, d[10], c1415, quotient[11], s1414, c1414);
addsub a14_15(s1316, d[09], c1416, quotient[11], s1415, c1415);
addsub a14_16(s1317, d[08], c1417, quotient[11], s1416, c1416);
addsub a14_17(s1318, d[07], c1418, quotient[11], s1417, c1417);
addsub a14_18(s1319, d[06], c1419, quotient[11], s1418, c1418);
addsub a14_19(s1320, d[05], c1420, quotient[11], s1419, c1419);
addsub a14_20(s1321, d[04], c1421, quotient[11], s1420, c1420);
addsub a14_21(s1322, d[03], c1422, quotient[11], s1421, c1421);
addsub a14_22(s1323, d[02], c1423, quotient[11], s1422, c1422);
addsub a14_23(s1324, d[01], c1424, quotient[11], s1423, c1423);
addsub a14_24(y[10], d[00], quotient[11], quotient[11], s1424, c1424);


addsub a15_00(s1401, d[24], c1501, quotient[10], s1500, quotient[09]);
addsub a15_01(s1402, d[23], c1502, quotient[10], s1501, c1501);
addsub a15_02(s1403, d[22], c1503, quotient[10], s1502, c1502);
addsub a15_03(s1404, d[21], c1504, quotient[10], s1503, c1503);
addsub a15_04(s1405, d[20], c1505, quotient[10], s1504, c1504);
addsub a15_05(s1406, d[19], c1506, quotient[10], s1505, c1505);
addsub a15_06(s1407, d[18], c1507, quotient[10], s1506, c1506);
addsub a15_07(s1408, d[17], c1508, quotient[10], s1507, c1507);
addsub a15_08(s1409, d[16], c1509, quotient[10], s1508, c1508);
addsub a15_09(s1410, d[15], c1510, quotient[10], s1509, c1509);
addsub a15_10(s1411, d[14], c1511, quotient[10], s1510, c1510);
addsub a15_11(s1412, d[13], c1512, quotient[10], s1511, c1511);
addsub a15_12(s1413, d[12], c1513, quotient[10], s1512, c1512);
addsub a15_13(s1414, d[11], c1514, quotient[10], s1513, c1513);
addsub a15_14(s1415, d[10], c1515, quotient[10], s1514, c1514);
addsub a15_15(s1416, d[09], c1516, quotient[10], s1515, c1515);
addsub a15_16(s1417, d[08], c1517, quotient[10], s1516, c1516);
addsub a15_17(s1418, d[07], c1518, quotient[10], s1517, c1517);
addsub a15_18(s1419, d[06], c1519, quotient[10], s1518, c1518);
addsub a15_19(s1420, d[05], c1520, quotient[10], s1519, c1519);
addsub a15_20(s1421, d[04], c1521, quotient[10], s1520, c1520);
addsub a15_21(s1422, d[03], c1522, quotient[10], s1521, c1521);
addsub a15_22(s1423, d[02], c1523, quotient[10], s1522, c1522);
addsub a15_23(s1424, d[01], c1524, quotient[10], s1523, c1523);
addsub a15_24(y[09], d[00], quotient[10], quotient[10], s1524, c1524);


addsub a16_00(s1501, d[24], c1601, quotient[09], s1600, quotient[08]);
addsub a16_01(s1502, d[23], c1602, quotient[09], s1601, c1601);
addsub a16_02(s1503, d[22], c1603, quotient[09], s1602, c1602);
addsub a16_03(s1504, d[21], c1604, quotient[09], s1603, c1603);
addsub a16_04(s1505, d[20], c1605, quotient[09], s1604, c1604);
addsub a16_05(s1506, d[19], c1606, quotient[09], s1605, c1605);
addsub a16_06(s1507, d[18], c1607, quotient[09], s1606, c1606);
addsub a16_07(s1508, d[17], c1608, quotient[09], s1607, c1607);
addsub a16_08(s1509, d[16], c1609, quotient[09], s1608, c1608);
addsub a16_09(s1510, d[15], c1610, quotient[09], s1609, c1609);
addsub a16_10(s1511, d[14], c1611, quotient[09], s1610, c1610);
addsub a16_11(s1512, d[13], c1612, quotient[09], s1611, c1611);
addsub a16_12(s1513, d[12], c1613, quotient[09], s1612, c1612);
addsub a16_13(s1514, d[11], c1614, quotient[09], s1613, c1613);
addsub a16_14(s1515, d[10], c1615, quotient[09], s1614, c1614);
addsub a16_15(s1516, d[09], c1616, quotient[09], s1615, c1615);
addsub a16_16(s1517, d[08], c1617, quotient[09], s1616, c1616);
addsub a16_17(s1518, d[07], c1618, quotient[09], s1617, c1617);
addsub a16_18(s1519, d[06], c1619, quotient[09], s1618, c1618);
addsub a16_19(s1520, d[05], c1620, quotient[09], s1619, c1619);
addsub a16_20(s1521, d[04], c1621, quotient[09], s1620, c1620);
addsub a16_21(s1522, d[03], c1622, quotient[09], s1621, c1621);
addsub a16_22(s1523, d[02], c1623, quotient[09], s1622, c1622);
addsub a16_23(s1524, d[01], c1624, quotient[09], s1623, c1623);
addsub a16_24(y[08], d[00], quotient[09], quotient[09], s1624, c1624);


addsub a17_00(s1601, d[24], c1701, quotient[08], s1700, quotient[07]);
addsub a17_01(s1602, d[23], c1702, quotient[08], s1701, c1701);
addsub a17_02(s1603, d[22], c1703, quotient[08], s1702, c1702);
addsub a17_03(s1604, d[21], c1704, quotient[08], s1703, c1703);
addsub a17_04(s1605, d[20], c1705, quotient[08], s1704, c1704);
addsub a17_05(s1606, d[19], c1706, quotient[08], s1705, c1705);
addsub a17_06(s1607, d[18], c1707, quotient[08], s1706, c1706);
addsub a17_07(s1608, d[17], c1708, quotient[08], s1707, c1707);
addsub a17_08(s1609, d[16], c1709, quotient[08], s1708, c1708);
addsub a17_09(s1610, d[15], c1710, quotient[08], s1709, c1709);
addsub a17_10(s1611, d[14], c1711, quotient[08], s1710, c1710);
addsub a17_11(s1612, d[13], c1712, quotient[08], s1711, c1711);
addsub a17_12(s1613, d[12], c1713, quotient[08], s1712, c1712);
addsub a17_13(s1614, d[11], c1714, quotient[08], s1713, c1713);
addsub a17_14(s1615, d[10], c1715, quotient[08], s1714, c1714);
addsub a17_15(s1616, d[09], c1716, quotient[08], s1715, c1715);
addsub a17_16(s1617, d[08], c1717, quotient[08], s1716, c1716);
addsub a17_17(s1618, d[07], c1718, quotient[08], s1717, c1717);
addsub a17_18(s1619, d[06], c1719, quotient[08], s1718, c1718);
addsub a17_19(s1620, d[05], c1720, quotient[08], s1719, c1719);
addsub a17_20(s1621, d[04], c1721, quotient[08], s1720, c1720);
addsub a17_21(s1622, d[03], c1722, quotient[08], s1721, c1721);
addsub a17_22(s1623, d[02], c1723, quotient[08], s1722, c1722);
addsub a17_23(s1624, d[01], c1724, quotient[08], s1723, c1723);
addsub a17_24(y[07], d[00], quotient[08], quotient[08], s1724, c1724);


addsub a18_00(s1701, d[24], c1801, quotient[07], s1800, quotient[06]);
addsub a18_01(s1702, d[23], c1802, quotient[07], s1801, c1801);
addsub a18_02(s1703, d[22], c1803, quotient[07], s1802, c1802);
addsub a18_03(s1704, d[21], c1804, quotient[07], s1803, c1803);
addsub a18_04(s1705, d[20], c1805, quotient[07], s1804, c1804);
addsub a18_05(s1706, d[19], c1806, quotient[07], s1805, c1805);
addsub a18_06(s1707, d[18], c1807, quotient[07], s1806, c1806);
addsub a18_07(s1708, d[17], c1808, quotient[07], s1807, c1807);
addsub a18_08(s1709, d[16], c1809, quotient[07], s1808, c1808);
addsub a18_09(s1710, d[15], c1810, quotient[07], s1809, c1809);
addsub a18_10(s1711, d[14], c1811, quotient[07], s1810, c1810);
addsub a18_11(s1712, d[13], c1812, quotient[07], s1811, c1811);
addsub a18_12(s1713, d[12], c1813, quotient[07], s1812, c1812);
addsub a18_13(s1714, d[11], c1814, quotient[07], s1813, c1813);
addsub a18_14(s1715, d[10], c1815, quotient[07], s1814, c1814);
addsub a18_15(s1716, d[09], c1816, quotient[07], s1815, c1815);
addsub a18_16(s1717, d[08], c1817, quotient[07], s1816, c1816);
addsub a18_17(s1718, d[07], c1818, quotient[07], s1817, c1817);
addsub a18_18(s1719, d[06], c1819, quotient[07], s1818, c1818);
addsub a18_19(s1720, d[05], c1820, quotient[07], s1819, c1819);
addsub a18_20(s1721, d[04], c1821, quotient[07], s1820, c1820);
addsub a18_21(s1722, d[03], c1822, quotient[07], s1821, c1821);
addsub a18_22(s1723, d[02], c1823, quotient[07], s1822, c1822);
addsub a18_23(s1724, d[01], c1824, quotient[07], s1823, c1823);
addsub a18_24(y[06], d[00], quotient[07], quotient[07], s1824, c1824);


addsub a19_00(s1801, d[24], c1901, quotient[06], s1900, quotient[05]);
addsub a19_01(s1802, d[23], c1902, quotient[06], s1901, c1901);
addsub a19_02(s1803, d[22], c1903, quotient[06], s1902, c1902);
addsub a19_03(s1804, d[21], c1904, quotient[06], s1903, c1903);
addsub a19_04(s1805, d[20], c1905, quotient[06], s1904, c1904);
addsub a19_05(s1806, d[19], c1906, quotient[06], s1905, c1905);
addsub a19_06(s1807, d[18], c1907, quotient[06], s1906, c1906);
addsub a19_07(s1808, d[17], c1908, quotient[06], s1907, c1907);
addsub a19_08(s1809, d[16], c1909, quotient[06], s1908, c1908);
addsub a19_09(s1810, d[15], c1910, quotient[06], s1909, c1909);
addsub a19_10(s1811, d[14], c1911, quotient[06], s1910, c1910);
addsub a19_11(s1812, d[13], c1912, quotient[06], s1911, c1911);
addsub a19_12(s1813, d[12], c1913, quotient[06], s1912, c1912);
addsub a19_13(s1814, d[11], c1914, quotient[06], s1913, c1913);
addsub a19_14(s1815, d[10], c1915, quotient[06], s1914, c1914);
addsub a19_15(s1816, d[09], c1916, quotient[06], s1915, c1915);
addsub a19_16(s1817, d[08], c1917, quotient[06], s1916, c1916);
addsub a19_17(s1818, d[07], c1918, quotient[06], s1917, c1917);
addsub a19_18(s1819, d[06], c1919, quotient[06], s1918, c1918);
addsub a19_19(s1820, d[05], c1920, quotient[06], s1919, c1919);
addsub a19_20(s1821, d[04], c1921, quotient[06], s1920, c1920);
addsub a19_21(s1822, d[03], c1922, quotient[06], s1921, c1921);
addsub a19_22(s1823, d[02], c1923, quotient[06], s1922, c1922);
addsub a19_23(s1824, d[01], c1924, quotient[06], s1923, c1923);
addsub a19_24(y[05], d[00], quotient[06], quotient[06], s1924, c1924);


addsub a20_00(s1901, d[24], c2001, quotient[05], s2000, quotient[04]);
addsub a20_01(s1902, d[23], c2002, quotient[05], s2001, c2001);
addsub a20_02(s1903, d[22], c2003, quotient[05], s2002, c2002);
addsub a20_03(s1904, d[21], c2004, quotient[05], s2003, c2003);
addsub a20_04(s1905, d[20], c2005, quotient[05], s2004, c2004);
addsub a20_05(s1906, d[19], c2006, quotient[05], s2005, c2005);
addsub a20_06(s1907, d[18], c2007, quotient[05], s2006, c2006);
addsub a20_07(s1908, d[17], c2008, quotient[05], s2007, c2007);
addsub a20_08(s1909, d[16], c2009, quotient[05], s2008, c2008);
addsub a20_09(s1910, d[15], c2010, quotient[05], s2009, c2009);
addsub a20_10(s1911, d[14], c2011, quotient[05], s2010, c2010);
addsub a20_11(s1912, d[13], c2012, quotient[05], s2011, c2011);
addsub a20_12(s1913, d[12], c2013, quotient[05], s2012, c2012);
addsub a20_13(s1914, d[11], c2014, quotient[05], s2013, c2013);
addsub a20_14(s1915, d[10], c2015, quotient[05], s2014, c2014);
addsub a20_15(s1916, d[09], c2016, quotient[05], s2015, c2015);
addsub a20_16(s1917, d[08], c2017, quotient[05], s2016, c2016);
addsub a20_17(s1918, d[07], c2018, quotient[05], s2017, c2017);
addsub a20_18(s1919, d[06], c2019, quotient[05], s2018, c2018);
addsub a20_19(s1920, d[05], c2020, quotient[05], s2019, c2019);
addsub a20_20(s1921, d[04], c2021, quotient[05], s2020, c2020);
addsub a20_21(s1922, d[03], c2022, quotient[05], s2021, c2021);
addsub a20_22(s1923, d[02], c2023, quotient[05], s2022, c2022);
addsub a20_23(s1924, d[01], c2024, quotient[05], s2023, c2023);
addsub a20_24(y[04], d[00], quotient[05], quotient[05], s2024, c2024);


addsub a21_00(s2001, d[24], c2101, quotient[04], s2100, quotient[03]);
addsub a21_01(s2002, d[23], c2102, quotient[04], s2101, c2101);
addsub a21_02(s2003, d[22], c2103, quotient[04], s2102, c2102);
addsub a21_03(s2004, d[21], c2104, quotient[04], s2103, c2103);
addsub a21_04(s2005, d[20], c2105, quotient[04], s2104, c2104);
addsub a21_05(s2006, d[19], c2106, quotient[04], s2105, c2105);
addsub a21_06(s2007, d[18], c2107, quotient[04], s2106, c2106);
addsub a21_07(s2008, d[17], c2108, quotient[04], s2107, c2107);
addsub a21_08(s2009, d[16], c2109, quotient[04], s2108, c2108);
addsub a21_09(s2010, d[15], c2110, quotient[04], s2109, c2109);
addsub a21_10(s2011, d[14], c2111, quotient[04], s2110, c2110);
addsub a21_11(s2012, d[13], c2112, quotient[04], s2111, c2111);
addsub a21_12(s2013, d[12], c2113, quotient[04], s2112, c2112);
addsub a21_13(s2014, d[11], c2114, quotient[04], s2113, c2113);
addsub a21_14(s2015, d[10], c2115, quotient[04], s2114, c2114);
addsub a21_15(s2016, d[09], c2116, quotient[04], s2115, c2115);
addsub a21_16(s2017, d[08], c2117, quotient[04], s2116, c2116);
addsub a21_17(s2018, d[07], c2118, quotient[04], s2117, c2117);
addsub a21_18(s2019, d[06], c2119, quotient[04], s2118, c2118);
addsub a21_19(s2020, d[05], c2120, quotient[04], s2119, c2119);
addsub a21_20(s2021, d[04], c2121, quotient[04], s2120, c2120);
addsub a21_21(s2022, d[03], c2122, quotient[04], s2121, c2121);
addsub a21_22(s2023, d[02], c2123, quotient[04], s2122, c2122);
addsub a21_23(s2024, d[01], c2124, quotient[04], s2123, c2123);
addsub a21_24(y[03], d[00], quotient[04], quotient[04], s2124, c2124);


addsub a22_00(s2101, d[24], c2201, quotient[03], s2200, quotient[02]);
addsub a22_01(s2102, d[23], c2202, quotient[03], s2201, c2201);
addsub a22_02(s2103, d[22], c2203, quotient[03], s2202, c2202);
addsub a22_03(s2104, d[21], c2204, quotient[03], s2203, c2203);
addsub a22_04(s2105, d[20], c2205, quotient[03], s2204, c2204);
addsub a22_05(s2106, d[19], c2206, quotient[03], s2205, c2205);
addsub a22_06(s2107, d[18], c2207, quotient[03], s2206, c2206);
addsub a22_07(s2108, d[17], c2208, quotient[03], s2207, c2207);
addsub a22_08(s2109, d[16], c2209, quotient[03], s2208, c2208);
addsub a22_09(s2110, d[15], c2210, quotient[03], s2209, c2209);
addsub a22_10(s2111, d[14], c2211, quotient[03], s2210, c2210);
addsub a22_11(s2112, d[13], c2212, quotient[03], s2211, c2211);
addsub a22_12(s2113, d[12], c2213, quotient[03], s2212, c2212);
addsub a22_13(s2114, d[11], c2214, quotient[03], s2213, c2213);
addsub a22_14(s2115, d[10], c2215, quotient[03], s2214, c2214);
addsub a22_15(s2116, d[09], c2216, quotient[03], s2215, c2215);
addsub a22_16(s2117, d[08], c2217, quotient[03], s2216, c2216);
addsub a22_17(s2118, d[07], c2218, quotient[03], s2217, c2217);
addsub a22_18(s2119, d[06], c2219, quotient[03], s2218, c2218);
addsub a22_19(s2120, d[05], c2220, quotient[03], s2219, c2219);
addsub a22_20(s2121, d[04], c2221, quotient[03], s2220, c2220);
addsub a22_21(s2122, d[03], c2222, quotient[03], s2221, c2221);
addsub a22_22(s2123, d[02], c2223, quotient[03], s2222, c2222);
addsub a22_23(s2124, d[01], c2224, quotient[03], s2223, c2223);
addsub a22_24(y[02], d[00], quotient[03], quotient[03], s2224, c2224);


addsub a23_00(s2201, d[24], c2301, quotient[02], s2300, quotient[01]);
addsub a23_01(s2202, d[23], c2302, quotient[02], s2301, c2301);
addsub a23_02(s2203, d[22], c2303, quotient[02], s2302, c2302);
addsub a23_03(s2204, d[21], c2304, quotient[02], s2303, c2303);
addsub a23_04(s2205, d[20], c2305, quotient[02], s2304, c2304);
addsub a23_05(s2206, d[19], c2306, quotient[02], s2305, c2305);
addsub a23_06(s2207, d[18], c2307, quotient[02], s2306, c2306);
addsub a23_07(s2208, d[17], c2308, quotient[02], s2307, c2307);
addsub a23_08(s2209, d[16], c2309, quotient[02], s2308, c2308);
addsub a23_09(s2210, d[15], c2310, quotient[02], s2309, c2309);
addsub a23_10(s2211, d[14], c2311, quotient[02], s2310, c2310);
addsub a23_11(s2212, d[13], c2312, quotient[02], s2311, c2311);
addsub a23_12(s2213, d[12], c2313, quotient[02], s2312, c2312);
addsub a23_13(s2214, d[11], c2314, quotient[02], s2313, c2313);
addsub a23_14(s2215, d[10], c2315, quotient[02], s2314, c2314);
addsub a23_15(s2216, d[09], c2316, quotient[02], s2315, c2315);
addsub a23_16(s2217, d[08], c2317, quotient[02], s2316, c2316);
addsub a23_17(s2218, d[07], c2318, quotient[02], s2317, c2317);
addsub a23_18(s2219, d[06], c2319, quotient[02], s2318, c2318);
addsub a23_19(s2220, d[05], c2320, quotient[02], s2319, c2319);
addsub a23_20(s2221, d[04], c2321, quotient[02], s2320, c2320);
addsub a23_21(s2222, d[03], c2322, quotient[02], s2321, c2321);
addsub a23_22(s2223, d[02], c2323, quotient[02], s2322, c2322);
addsub a23_23(s2224, d[01], c2324, quotient[02], s2323, c2323);
addsub a23_24(y[01], d[00], quotient[02], quotient[02], s2324, c2324);


addsub a24_00(s2301, d[24], c2401, quotient[01], s2400, quotient[00]);
addsub a24_01(s2302, d[23], c2402, quotient[01], s2401, c2401);
addsub a24_02(s2303, d[22], c2403, quotient[01], s2402, c2402);
addsub a24_03(s2304, d[21], c2404, quotient[01], s2403, c2403);
addsub a24_04(s2305, d[20], c2405, quotient[01], s2404, c2404);
addsub a24_05(s2306, d[19], c2406, quotient[01], s2405, c2405);
addsub a24_06(s2307, d[18], c2407, quotient[01], s2406, c2406);
addsub a24_07(s2308, d[17], c2408, quotient[01], s2407, c2407);
addsub a24_08(s2309, d[16], c2409, quotient[01], s2408, c2408);
addsub a24_09(s2310, d[15], c2410, quotient[01], s2409, c2409);
addsub a24_10(s2311, d[14], c2411, quotient[01], s2410, c2410);
addsub a24_11(s2312, d[13], c2412, quotient[01], s2411, c2411);
addsub a24_12(s2313, d[12], c2413, quotient[01], s2412, c2412);
addsub a24_13(s2314, d[11], c2414, quotient[01], s2413, c2413);
addsub a24_14(s2315, d[10], c2415, quotient[01], s2414, c2414);
addsub a24_15(s2316, d[09], c2416, quotient[01], s2415, c2415);
addsub a24_16(s2317, d[08], c2417, quotient[01], s2416, c2416);
addsub a24_17(s2318, d[07], c2418, quotient[01], s2417, c2417);
addsub a24_18(s2319, d[06], c2419, quotient[01], s2418, c2418);
addsub a24_19(s2320, d[05], c2420, quotient[01], s2419, c2419);
addsub a24_20(s2321, d[04], c2421, quotient[01], s2420, c2420);
addsub a24_21(s2322, d[03], c2422, quotient[01], s2421, c2421);
addsub a24_22(s2323, d[02], c2423, quotient[01], s2422, c2422);
addsub a24_23(s2324, d[01], c2424, quotient[01], s2423, c2423);
addsub a24_24(y[00], d[00], quotient[01], quotient[01], s2424, c2424);


assign remainder = s2400 ? {s2400,s2401,s2402,s2403,s2404,s2405,s2406,s2407,s2408,s2409,s2410,s2411,s2412,s2413,s2414,s2415,s2416,s2417,s2418,s2419,s2420,s2421,s2422,s2423,s2424} + divisor : {s2400,s2401,s2402,s2403,s2404,s2405,s2406,s2407,s2408,s2409,s2410,s2411,s2412,s2413,s2414,s2415,s2416,s2417,s2418,s2419,s2420,s2421,s2422,s2423,s2424};

always @(posedge clk) begin
    if (rst) begin
        y <= { 24'b0, dividend };
        d <= { 1'b0, divisor };
    end
end
endmodule
